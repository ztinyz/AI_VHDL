library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package weights_pkg is
  type conv1_weight_32_1_3_3_t is array (0 to 287) of std_logic_vector(7 downto 0);
  constant conv1_weight : conv1_weight_32_1_3_3_t := (
    x"1b", x"36", x"0f", x"d4", x"c2", x"08", x"e8", x"f7",
    x"d3", x"e3", x"18", x"fe", x"a4", x"18", x"21", x"65",
    x"82", x"df", x"0e", x"01", x"06", x"92", x"83", x"d7",
    x"8d", x"f2", x"50", x"eb", x"1c", x"e4", x"25", x"f2",
    x"cd", x"a9", x"f3", x"03", x"f7", x"24", x"0b", x"04",
    x"1c", x"14", x"ea", x"30", x"ff", x"dc", x"ee", x"32",
    x"f9", x"30", x"f7", x"28", x"f8", x"dc", x"d0", x"c9",
    x"d5", x"04", x"f4", x"e1", x"18", x"1f", x"24", x"03",
    x"1d", x"ff", x"ee", x"d7", x"eb", x"04", x"ea", x"f3",
    x"00", x"df", x"1e", x"fc", x"3d", x"87", x"06", x"00",
    x"36", x"f4", x"df", x"f1", x"e8", x"ee", x"00", x"0b",
    x"f9", x"03", x"09", x"fd", x"4b", x"f4", x"8e", x"f5",
    x"36", x"f8", x"10", x"ff", x"54", x"04", x"fa", x"d5",
    x"28", x"db", x"0b", x"19", x"0b", x"e0", x"e7", x"28",
    x"7a", x"e6", x"da", x"58", x"0a", x"03", x"fe", x"d1",
    x"da", x"36", x"bf", x"89", x"0f", x"f9", x"0a", x"0c",
    x"0c", x"fe", x"00", x"f5", x"54", x"a1", x"23", x"4d",
    x"f2", x"b3", x"eb", x"90", x"93", x"91", x"91", x"b9",
    x"09", x"01", x"d9", x"05", x"a7", x"54", x"0a", x"0f",
    x"02", x"f9", x"f3", x"17", x"e4", x"fb", x"16", x"ea",
    x"36", x"02", x"df", x"e6", x"f6", x"20", x"26", x"14",
    x"e4", x"b5", x"db", x"13", x"fb", x"f4", x"23", x"fe",
    x"40", x"1f", x"22", x"fe", x"22", x"f8", x"c8", x"ef",
    x"d1", x"fd", x"e9", x"4d", x"03", x"fa", x"d2", x"c4",
    x"06", x"15", x"7a", x"14", x"22", x"c9", x"24", x"d1",
    x"eb", x"28", x"e0", x"fc", x"1a", x"f0", x"00", x"1e",
    x"0a", x"23", x"26", x"e1", x"84", x"f1", x"46", x"b5",
    x"a6", x"e7", x"ef", x"a2", x"5c", x"9d", x"d8", x"ef",
    x"dc", x"16", x"e8", x"d1", x"0c", x"53", x"0d", x"e9",
    x"f4", x"1e", x"f2", x"f6", x"19", x"d9", x"ed", x"21",
    x"ce", x"e8", x"12", x"13", x"2a", x"04", x"26", x"07",
    x"42", x"0c", x"d5", x"ed", x"f8", x"2e", x"de", x"1a",
    x"0b", x"dc", x"1d", x"ff", x"f2", x"ff", x"e7", x"40",
    x"04", x"fe", x"dd", x"dd", x"b3", x"fd", x"eb", x"f2",
    x"eb", x"a1", x"04", x"c6", x"a2", x"fa", x"c4", x"10",
    x"11", x"13", x"15", x"16", x"f6", x"d6", x"af", x"73"
  );

  type conv1_bias_32_t is array (0 to 31) of std_logic_vector(7 downto 0);
  constant conv1_bias : conv1_bias_32_t := (
    x"e1", x"fb", x"d3", x"fc", x"b3", x"cb", x"f0", x"db",
    x"c2", x"ee", x"be", x"ac", x"fe", x"f8", x"b4", x"e2",
    x"c6", x"d5", x"fe", x"9b", x"d2", x"ff", x"e1", x"ae",
    x"f0", x"c1", x"f3", x"9f", x"da", x"f9", x"1e", x"e8"
  );

  type conv1_activation_post_process_eps_1_t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant conv1_activation_post_process_eps : conv1_activation_post_process_eps_1_t := (
    x"00"
  );

  type conv1_activation_post_process_min_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant conv1_activation_post_process_min_val : conv1_activation_post_process_min_val__t := (
    x"9b"
  );

  type conv1_activation_post_process_max_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant conv1_activation_post_process_max_val : conv1_activation_post_process_max_val__t := (
    x"1e"
  );

  type conv2_weight_64_32_3_3_t is array (0 to 18431) of std_logic_vector(7 downto 0);
  constant conv2_weight : conv2_weight_64_32_3_3_t := (
    x"24", x"e4", x"bb", x"a0", x"af", x"66", x"f2", x"ef",
    x"b9", x"09", x"eb", x"fb", x"2c", x"d3", x"aa", x"3e",
    x"d4", x"dc", x"be", x"07", x"fb", x"16", x"09", x"fd",
    x"e4", x"05", x"b6", x"f4", x"aa", x"01", x"d3", x"10",
    x"20", x"72", x"35", x"fb", x"ee", x"e0", x"1f", x"d2",
    x"d7", x"54", x"86", x"10", x"45", x"32", x"de", x"de",
    x"c7", x"e9", x"e0", x"2c", x"1f", x"0a", x"55", x"ff",
    x"1f", x"f3", x"04", x"df", x"9d", x"d3", x"fd", x"fe",
    x"fd", x"03", x"00", x"05", x"ff", x"fe", x"05", x"03",
    x"13", x"e8", x"21", x"f4", x"c3", x"d5", x"35", x"b5",
    x"c6", x"f9", x"ff", x"fb", x"fa", x"00", x"06", x"07",
    x"ff", x"01", x"e8", x"02", x"43", x"d1", x"34", x"00",
    x"b1", x"28", x"ea", x"5a", x"01", x"03", x"e6", x"fd",
    x"1b", x"d9", x"f6", x"25", x"c4", x"dc", x"f5", x"cf",
    x"f7", x"07", x"d0", x"12", x"12", x"fe", x"e9", x"02",
    x"f6", x"00", x"fa", x"af", x"ec", x"04", x"f3", x"47",
    x"fc", x"64", x"38", x"d2", x"8d", x"0a", x"e0", x"f8",
    x"96", x"28", x"b9", x"55", x"37", x"ab", x"09", x"fd",
    x"9e", x"d3", x"01", x"fe", x"09", x"00", x"da", x"14",
    x"e9", x"d5", x"d4", x"26", x"ff", x"ec", x"2b", x"b1",
    x"25", x"2a", x"bc", x"cc", x"1d", x"d0", x"dd", x"17",
    x"06", x"fc", x"0b", x"e9", x"e6", x"dc", x"5a", x"09",
    x"23", x"a8", x"a4", x"fd", x"bc", x"d9", x"be", x"af",
    x"b3", x"d2", x"c3", x"c0", x"04", x"70", x"fe", x"10",
    x"81", x"94", x"0b", x"87", x"08", x"2f", x"d5", x"ff",
    x"20", x"85", x"ec", x"12", x"2f", x"8a", x"0b", x"f5",
    x"eb", x"fb", x"bf", x"fa", x"27", x"82", x"e9", x"0b",
    x"2a", x"8e", x"29", x"ee", x"ec", x"16", x"31", x"f7",
    x"fa", x"ab", x"cc", x"14", x"c8", x"ea", x"09", x"bb",
    x"e2", x"df", x"d4", x"12", x"13", x"fb", x"14", x"11",
    x"df", x"18", x"3b", x"24", x"d0", x"f8", x"94", x"bc",
    x"2f", x"b8", x"f5", x"02", x"2d", x"b6", x"36", x"ec",
    x"ae", x"fa", x"86", x"e9", x"32", x"f7", x"e7", x"fb",
    x"c2", x"f6", x"05", x"1c", x"e9", x"12", x"f1", x"f3",
    x"e0", x"00", x"05", x"ee", x"fe", x"e8", x"ba", x"16",
    x"c8", x"e8", x"a9", x"8d", x"d8", x"f1", x"dd", x"fa",
    x"1d", x"04", x"3c", x"01", x"f8", x"26", x"19", x"e8",
    x"e4", x"12", x"0a", x"04", x"25", x"3e", x"29", x"33",
    x"4f", x"02", x"3a", x"12", x"1c", x"f0", x"de", x"51",
    x"15", x"51", x"8d", x"17", x"16", x"06", x"1b", x"1a",
    x"fd", x"1a", x"09", x"46", x"d9", x"f9", x"19", x"e6",
    x"9d", x"bb", x"04", x"f0", x"cb", x"27", x"fd", x"e9",
    x"01", x"d4", x"aa", x"14", x"9b", x"66", x"2b", x"05",
    x"3f", x"1a", x"e6", x"c9", x"2f", x"2a", x"d0", x"02",
    x"06", x"fa", x"04", x"02", x"f9", x"f9", x"ff", x"fa",
    x"14", x"16", x"99", x"1a", x"12", x"76", x"cb", x"db",
    x"23", x"fa", x"04", x"f9", x"f9", x"fb", x"fd", x"03",
    x"02", x"f9", x"24", x"4a", x"12", x"0b", x"12", x"14",
    x"1a", x"0b", x"e4", x"fa", x"25", x"f8", x"fe", x"ec",
    x"ef", x"12", x"23", x"61", x"20", x"0b", x"ec", x"2f",
    x"00", x"bb", x"20", x"49", x"28", x"fa", x"d9", x"21",
    x"02", x"02", x"b9", x"18", x"2a", x"42", x"ea", x"11",
    x"0c", x"00", x"0d", x"df", x"fb", x"2d", x"ef", x"38",
    x"39", x"0b", x"22", x"07", x"0b", x"ee", x"07", x"d3",
    x"2d", x"de", x"53", x"12", x"c3", x"2a", x"09", x"0f",
    x"b2", x"fd", x"02", x"f2", x"e8", x"7f", x"55", x"e4",
    x"fc", x"80", x"fb", x"da", x"18", x"fd", x"dc", x"d6",
    x"19", x"25", x"cd", x"13", x"19", x"46", x"12", x"e9",
    x"c2", x"06", x"f1", x"b3", x"f0", x"c8", x"dc", x"e6",
    x"06", x"e4", x"37", x"07", x"19", x"e9", x"bb", x"db",
    x"1d", x"fb", x"e6", x"19", x"1c", x"3b", x"f9", x"f0",
    x"d5", x"35", x"ff", x"d8", x"f5", x"03", x"18", x"de",
    x"e4", x"16", x"1f", x"28", x"38", x"18", x"06", x"34",
    x"2f", x"20", x"0d", x"f9", x"df", x"c1", x"f7", x"29",
    x"01", x"de", x"d7", x"1b", x"24", x"19", x"c4", x"ec",
    x"2b", x"e6", x"04", x"07", x"28", x"aa", x"ea", x"e0",
    x"ef", x"f9", x"c9", x"e3", x"f7", x"32", x"1b", x"16",
    x"0f", x"f8", x"17", x"05", x"12", x"09", x"e8", x"29",
    x"00", x"cf", x"d5", x"d6", x"e0", x"ec", x"0b", x"45",
    x"e9", x"e0", x"ef", x"26", x"37", x"d8", x"1f", x"e4",
    x"df", x"ef", x"f8", x"e6", x"b7", x"ee", x"ee", x"21",
    x"0b", x"1f", x"1b", x"ba", x"fe", x"19", x"1b", x"e6",
    x"e9", x"24", x"54", x"f5", x"05", x"16", x"d6", x"03",
    x"08", x"1a", x"09", x"32", x"69", x"28", x"31", x"c2",
    x"24", x"27", x"dd", x"05", x"03", x"e2", x"0e", x"23",
    x"37", x"f8", x"25", x"04", x"30", x"29", x"f2", x"f3",
    x"e2", x"e9", x"0f", x"a4", x"ee", x"df", x"2e", x"ea",
    x"fe", x"33", x"f2", x"18", x"1b", x"e6", x"19", x"ca",
    x"b4", x"f7", x"12", x"3e", x"26", x"d0", x"21", x"03",
    x"08", x"f0", x"07", x"d4", x"cc", x"29", x"e3", x"fa",
    x"fa", x"fc", x"fb", x"02", x"04", x"06", x"05", x"fb",
    x"06", x"0e", x"01", x"05", x"07", x"fa", x"3e", x"22",
    x"ff", x"fd", x"fd", x"03", x"02", x"00", x"fc", x"fb",
    x"01", x"06", x"03", x"26", x"06", x"e0", x"58", x"07",
    x"3d", x"04", x"22", x"81", x"f0", x"00", x"f7", x"34",
    x"17", x"0e", x"ff", x"15", x"58", x"0e", x"f5", x"bf",
    x"fe", x"1f", x"fb", x"e2", x"f8", x"1a", x"2c", x"0f",
    x"0c", x"f7", x"01", x"75", x"c6", x"f6", x"c7", x"1f",
    x"11", x"ef", x"d7", x"dc", x"26", x"ff", x"08", x"ec",
    x"44", x"27", x"f8", x"9d", x"1a", x"53", x"ad", x"b0",
    x"ff", x"0a", x"dd", x"e9", x"1a", x"24", x"3d", x"35",
    x"0b", x"0f", x"fc", x"f2", x"0b", x"0b", x"5c", x"11",
    x"ed", x"ec", x"ff", x"2b", x"3c", x"38", x"21", x"b5",
    x"0c", x"10", x"e7", x"bb", x"08", x"f5", x"dc", x"f2",
    x"28", x"f3", x"18", x"fb", x"1d", x"4a", x"0e", x"10",
    x"26", x"d7", x"2d", x"17", x"14", x"d3", x"01", x"1a",
    x"99", x"a7", x"18", x"bb", x"17", x"39", x"b8", x"bd",
    x"13", x"fe", x"c3", x"ed", x"39", x"3c", x"47", x"fe",
    x"e9", x"1b", x"ff", x"c8", x"02", x"d4", x"35", x"4b",
    x"2b", x"19", x"19", x"18", x"04", x"41", x"07", x"41",
    x"d2", x"da", x"1a", x"f0", x"10", x"fe", x"ff", x"0d",
    x"38", x"fc", x"fb", x"f9", x"21", x"ec", x"db", x"31",
    x"f6", x"d8", x"cd", x"dd", x"e9", x"e9", x"d1", x"e5",
    x"0e", x"06", x"15", x"44", x"14", x"f2", x"ef", x"aa",
    x"62", x"19", x"a3", x"1b", x"24", x"f1", x"2f", x"49",
    x"36", x"16", x"e9", x"03", x"e9", x"cc", x"10", x"dc",
    x"bf", x"ee", x"0e", x"aa", x"e8", x"b6", x"84", x"00",
    x"0a", x"fd", x"18", x"dc", x"f2", x"2a", x"e8", x"f2",
    x"e9", x"f2", x"ed", x"80", x"77", x"e6", x"ae", x"7c",
    x"d1", x"96", x"f3", x"03", x"20", x"e4", x"ef", x"1a",
    x"c6", x"e7", x"37", x"d3", x"f4", x"ff", x"dc", x"d7",
    x"34", x"53", x"88", x"aa", x"01", x"f5", x"38", x"e6",
    x"d3", x"bc", x"fa", x"d0", x"a8", x"d9", x"ef", x"08",
    x"06", x"d5", x"06", x"2a", x"bf", x"ca", x"d2", x"ce",
    x"f6", x"fc", x"c5", x"e8", x"3f", x"ee", x"22", x"fc",
    x"32", x"f1", x"f2", x"ff", x"74", x"e7", x"d8", x"04",
    x"fa", x"fc", x"fe", x"fd", x"00", x"fa", x"05", x"f9",
    x"b7", x"cd", x"eb", x"04", x"f7", x"ac", x"f3", x"0c",
    x"dc", x"03", x"fa", x"fe", x"fa", x"ff", x"07", x"fb",
    x"03", x"fb", x"22", x"11", x"35", x"dd", x"0f", x"11",
    x"87", x"0c", x"fd", x"9e", x"ee", x"28", x"d1", x"6e",
    x"20", x"fb", x"a4", x"f6", x"a2", x"d8", x"c8", x"a3",
    x"e1", x"ec", x"9d", x"bc", x"83", x"c9", x"60", x"1b",
    x"08", x"71", x"14", x"09", x"eb", x"d2", x"c6", x"a8",
    x"dd", x"d3", x"03", x"a9", x"fc", x"04", x"f3", x"cc",
    x"eb", x"b4", x"bb", x"c8", x"bf", x"a1", x"f4", x"99",
    x"93", x"ff", x"ec", x"e2", x"b2", x"f0", x"7b", x"bc",
    x"ce", x"c8", x"93", x"04", x"18", x"7a", x"d1", x"fd",
    x"07", x"bf", x"01", x"d7", x"11", x"ea", x"fa", x"d0",
    x"dc", x"1d", x"a5", x"27", x"e4", x"f3", x"43", x"19",
    x"dd", x"45", x"36", x"fc", x"ee", x"c3", x"1e", x"1b",
    x"e1", x"a4", x"10", x"33", x"e5", x"0b", x"fd", x"f7",
    x"10", x"0d", x"ce", x"fd", x"10", x"00", x"cd", x"e2",
    x"cd", x"f8", x"ee", x"bd", x"ce", x"05", x"d1", x"e9",
    x"cf", x"0e", x"8a", x"16", x"c2", x"25", x"5f", x"cf",
    x"7d", x"c4", x"01", x"89", x"b2", x"ef", x"93", x"ab",
    x"e7", x"2d", x"a5", x"1f", x"11", x"e8", x"f2", x"02",
    x"11", x"b3", x"0d", x"f2", x"12", x"ce", x"06", x"ed",
    x"d6", x"a7", x"e2", x"a9", x"af", x"f0", x"f4", x"e6",
    x"b2", x"eb", x"d6", x"95", x"02", x"db", x"f9", x"00",
    x"0a", x"dd", x"02", x"07", x"b6", x"e5", x"0b", x"27",
    x"98", x"b7", x"1e", x"7d", x"9a", x"ee", x"54", x"ff",
    x"10", x"26", x"f6", x"03", x"2c", x"f9", x"ff", x"f8",
    x"ff", x"ed", x"d5", x"aa", x"0e", x"db", x"a9", x"93",
    x"6d", x"dc", x"cb", x"67", x"84", x"0a", x"9b", x"f7",
    x"05", x"3c", x"11", x"bd", x"f9", x"d5", x"fa", x"f6",
    x"18", x"09", x"5a", x"94", x"c7", x"31", x"44", x"0e",
    x"02", x"0d", x"5a", x"26", x"27", x"c0", x"bc", x"f8",
    x"06", x"ff", x"19", x"f1", x"f8", x"ed", x"03", x"04",
    x"38", x"09", x"20", x"ee", x"f4", x"32", x"e4", x"03",
    x"16", x"26", x"2e", x"36", x"09", x"03", x"1c", x"e5",
    x"d6", x"0f", x"0c", x"f7", x"b2", x"95", x"0c", x"06",
    x"07", x"02", x"04", x"fe", x"00", x"fd", x"07", x"07",
    x"18", x"f0", x"1c", x"06", x"f1", x"da", x"2a", x"61",
    x"06", x"05", x"fa", x"00", x"fe", x"06", x"fd", x"06",
    x"03", x"fe", x"16", x"19", x"02", x"1a", x"c8", x"f6",
    x"e4", x"11", x"28", x"f5", x"1d", x"fc", x"4c", x"38",
    x"14", x"ce", x"e5", x"0e", x"2c", x"c5", x"82", x"e1",
    x"e8", x"ee", x"0d", x"12", x"08", x"16", x"db", x"ae",
    x"e0", x"e3", x"09", x"2c", x"41", x"0e", x"13", x"0c",
    x"04", x"cf", x"32", x"22", x"47", x"0c", x"04", x"f8",
    x"b4", x"c8", x"a1", x"7e", x"ec", x"0d", x"39", x"65",
    x"fe", x"db", x"27", x"f2", x"00", x"1d", x"fd", x"1b",
    x"43", x"06", x"d6", x"e9", x"fb", x"30", x"1e", x"02",
    x"ff", x"fe", x"20", x"c7", x"ba", x"e2", x"f9", x"1d",
    x"e9", x"fe", x"22", x"f0", x"02", x"1c", x"29", x"04",
    x"0d", x"b3", x"ee", x"3a", x"17", x"0f", x"13", x"da",
    x"e4", x"f0", x"91", x"40", x"1b", x"ee", x"af", x"db",
    x"b1", x"e8", x"13", x"82", x"04", x"3d", x"42", x"19",
    x"16", x"dc", x"c8", x"f1", x"10", x"17", x"d5", x"2a",
    x"fe", x"0c", x"ac", x"d5", x"3c", x"01", x"e9", x"fd",
    x"4f", x"0c", x"18", x"ac", x"4d", x"fa", x"44", x"45",
    x"1b", x"0f", x"00", x"fa", x"0d", x"05", x"37", x"79",
    x"ed", x"fc", x"12", x"b7", x"15", x"f3", x"1c", x"d6",
    x"37", x"f7", x"21", x"41", x"16", x"f5", x"05", x"f6",
    x"17", x"ec", x"2c", x"e6", x"6c", x"ea", x"2b", x"ec",
    x"05", x"01", x"33", x"ca", x"eb", x"3f", x"3f", x"e5",
    x"1d", x"dc", x"20", x"aa", x"1d", x"0c", x"d3", x"cb",
    x"ee", x"08", x"08", x"a4", x"03", x"e8", x"cd", x"13",
    x"9a", x"b9", x"e1", x"d0", x"f7", x"f9", x"d7", x"ef",
    x"e8", x"af", x"d9", x"09", x"22", x"51", x"0a", x"2f",
    x"27", x"03", x"b9", x"9c", x"ca", x"f1", x"2d", x"d3",
    x"23", x"28", x"00", x"d9", x"ef", x"f1", x"0c", x"50",
    x"72", x"48", x"3d", x"09", x"0b", x"20", x"1f", x"1f",
    x"21", x"1c", x"1f", x"31", x"0b", x"03", x"1d", x"15",
    x"da", x"a3", x"24", x"9a", x"6d", x"00", x"31", x"36",
    x"06", x"f9", x"d9", x"e8", x"71", x"8a", x"fa", x"aa",
    x"d9", x"12", x"e7", x"0e", x"24", x"24", x"fa", x"fd",
    x"fb", x"06", x"02", x"07", x"07", x"05", x"fd", x"02",
    x"11", x"10", x"0b", x"16", x"fc", x"b4", x"d2", x"dc",
    x"9b", x"01", x"f9", x"05", x"05", x"06", x"03", x"06",
    x"ff", x"05", x"15", x"ed", x"65", x"05", x"a4", x"a6",
    x"28", x"0c", x"dc", x"2b", x"12", x"47", x"da", x"0c",
    x"ad", x"fc", x"f8", x"c7", x"fe", x"10", x"f8", x"0b",
    x"18", x"d9", x"fa", x"f6", x"f0", x"0a", x"bf", x"74",
    x"e7", x"08", x"44", x"1b", x"23", x"d6", x"15", x"0a",
    x"01", x"f0", x"e9", x"af", x"27", x"01", x"79", x"1b",
    x"ee", x"fd", x"0a", x"b4", x"de", x"4c", x"35", x"54",
    x"1d", x"1e", x"81", x"ea", x"f9", x"00", x"f0", x"d6",
    x"f9", x"1c", x"1a", x"ba", x"04", x"c0", x"d2", x"07",
    x"11", x"47", x"fd", x"c8", x"e0", x"17", x"27", x"4c",
    x"1a", x"16", x"64", x"f5", x"0a", x"e9", x"02", x"36",
    x"47", x"0e", x"14", x"32", x"e7", x"21", x"59", x"dd",
    x"48", x"6e", x"f6", x"fb", x"5b", x"19", x"0f", x"cd",
    x"13", x"4a", x"43", x"e6", x"b2", x"ff", x"16", x"1e",
    x"17", x"13", x"fb", x"d5", x"f8", x"fe", x"cb", x"e9",
    x"03", x"06", x"de", x"02", x"fb", x"1f", x"30", x"c7",
    x"28", x"66", x"21", x"16", x"f5", x"00", x"f9", x"ea",
    x"0a", x"15", x"f4", x"a4", x"d7", x"24", x"1f", x"0d",
    x"13", x"23", x"ee", x"d3", x"11", x"c8", x"dd", x"98",
    x"00", x"df", x"43", x"cf", x"ec", x"75", x"14", x"34",
    x"00", x"08", x"2a", x"27", x"07", x"23", x"23", x"04",
    x"de", x"a9", x"10", x"e0", x"af", x"e7", x"07", x"b5",
    x"e0", x"0d", x"51", x"e8", x"08", x"49", x"d3", x"f3",
    x"df", x"c9", x"ec", x"e7", x"c4", x"ea", x"d9", x"07",
    x"ca", x"da", x"2b", x"0c", x"04", x"0c", x"07", x"4a",
    x"d8", x"f1", x"cb", x"ee", x"0a", x"ca", x"cd", x"03",
    x"d1", x"1a", x"ed", x"f1", x"0c", x"f4", x"81", x"57",
    x"1d", x"25", x"de", x"17", x"0a", x"38", x"17", x"f4",
    x"4c", x"f8", x"e4", x"00", x"bd", x"fd", x"a7", x"0f",
    x"20", x"07", x"18", x"00", x"1a", x"07", x"16", x"a7",
    x"00", x"f5", x"fa", x"d7", x"c5", x"0e", x"f5", x"1e",
    x"06", x"07", x"09", x"07", x"e9", x"32", x"02", x"03",
    x"cc", x"d6", x"ca", x"c1", x"ed", x"e2", x"b1", x"05",
    x"07", x"06", x"ff", x"04", x"fc", x"03", x"01", x"01",
    x"09", x"cd", x"e0", x"ca", x"05", x"36", x"ff", x"f3",
    x"1b", x"fc", x"f9", x"01", x"fb", x"ff", x"05", x"05",
    x"fc", x"fe", x"08", x"bb", x"ca", x"e7", x"ef", x"c3",
    x"c8", x"93", x"0f", x"eb", x"09", x"04", x"03", x"ff",
    x"de", x"73", x"7e", x"c8", x"f8", x"f2", x"2c", x"2f",
    x"2f", x"07", x"3b", x"36", x"f3", x"ec", x"0d", x"c3",
    x"a7", x"f7", x"b7", x"dd", x"02", x"da", x"f6", x"da",
    x"08", x"d2", x"f2", x"07", x"d0", x"08", x"62", x"1f",
    x"ef", x"45", x"e6", x"18", x"21", x"eb", x"42", x"0c",
    x"eb", x"15", x"0b", x"ee", x"30", x"1e", x"24", x"e2",
    x"0b", x"df", x"09", x"1b", x"0b", x"23", x"e1", x"28",
    x"3f", x"57", x"e6", x"04", x"f2", x"ff", x"25", x"10",
    x"f8", x"2a", x"d1", x"33", x"f5", x"16", x"d2", x"df",
    x"d1", x"44", x"ed", x"c1", x"09", x"d1", x"0f", x"1d",
    x"f1", x"17", x"22", x"04", x"0d", x"82", x"e2", x"ac",
    x"df", x"f5", x"c5", x"0e", x"fa", x"d2", x"e7", x"dd",
    x"fd", x"83", x"0c", x"0c", x"64", x"f1", x"c1", x"13",
    x"1d", x"e9", x"05", x"da", x"c7", x"1d", x"b1", x"9f",
    x"1a", x"12", x"1d", x"f2", x"2e", x"22", x"4b", x"18",
    x"ff", x"f1", x"0b", x"d8", x"89", x"b0", x"95", x"5d",
    x"a4", x"8c", x"e2", x"01", x"10", x"dc", x"05", x"eb",
    x"4d", x"15", x"a9", x"b6", x"f4", x"03", x"90", x"dd",
    x"06", x"9d", x"8f", x"ee", x"00", x"24", x"0a", x"be",
    x"18", x"11", x"1b", x"16", x"d2", x"18", x"cd", x"19",
    x"e8", x"f4", x"ef", x"f8", x"2c", x"a4", x"eb", x"15",
    x"f2", x"0d", x"25", x"ec", x"2c", x"14", x"d6", x"ea",
    x"b4", x"f6", x"e3", x"a4", x"d7", x"2d", x"1b", x"d8",
    x"04", x"9a", x"09", x"0a", x"2a", x"27", x"fd", x"18",
    x"42", x"e9", x"b6", x"0d", x"fa", x"f8", x"0d", x"00",
    x"2f", x"02", x"de", x"1b", x"f1", x"bf", x"d8", x"dd",
    x"06", x"1b", x"15", x"de", x"10", x"46", x"df", x"16",
    x"da", x"db", x"b8", x"ec", x"15", x"2c", x"00", x"f6",
    x"09", x"17", x"e7", x"d0", x"ef", x"03", x"2a", x"31",
    x"1f", x"04", x"e0", x"0b", x"9d", x"ef", x"d3", x"c4",
    x"f1", x"df", x"cc", x"f3", x"b0", x"de", x"03", x"fa",
    x"07", x"00", x"fe", x"04", x"04", x"07", x"01", x"fe",
    x"26", x"08", x"02", x"44", x"0d", x"0c", x"cc", x"80",
    x"d8", x"ff", x"07", x"05", x"03", x"ff", x"fe", x"04",
    x"fe", x"fe", x"12", x"e8", x"0f", x"c4", x"d4", x"20",
    x"fb", x"18", x"29", x"37", x"d8", x"0f", x"34", x"0b",
    x"f1", x"af", x"3b", x"26", x"b1", x"11", x"37", x"2c",
    x"9f", x"e6", x"ca", x"c6", x"be", x"4f", x"34", x"d6",
    x"3d", x"42", x"0e", x"b4", x"01", x"f3", x"1c", x"f4",
    x"1e", x"02", x"16", x"1e", x"8a", x"ee", x"17", x"d4",
    x"d3", x"fb", x"24", x"8f", x"8e", x"26", x"c8", x"b5",
    x"ee", x"23", x"1a", x"21", x"0a", x"13", x"8f", x"af",
    x"c3", x"d1", x"33", x"13", x"f5", x"0b", x"c5", x"01",
    x"ea", x"d4", x"09", x"bb", x"23", x"e3", x"ce", x"48",
    x"13", x"9a", x"0f", x"30", x"d6", x"21", x"db", x"fd",
    x"34", x"ad", x"33", x"e9", x"d0", x"f0", x"3b", x"ef",
    x"0c", x"1f", x"b4", x"de", x"b2", x"07", x"ff", x"de",
    x"d8", x"28", x"bb", x"12", x"00", x"cb", x"45", x"6b",
    x"fb", x"05", x"f6", x"e8", x"5d", x"7b", x"b2", x"7b",
    x"69", x"de", x"37", x"25", x"dd", x"ec", x"f1", x"ff",
    x"dd", x"f1", x"4a", x"b9", x"f1", x"63", x"02", x"a8",
    x"19", x"07", x"e8", x"f2", x"cd", x"04", x"14", x"36",
    x"03", x"26", x"ef", x"50", x"f3", x"07", x"1b", x"e0",
    x"fa", x"e1", x"e7", x"d4", x"c2", x"fe", x"02", x"28",
    x"fb", x"ef", x"3a", x"e7", x"37", x"5e", x"01", x"d2",
    x"ef", x"08", x"9f", x"51", x"de", x"b4", x"ee", x"2f",
    x"1f", x"06", x"21", x"12", x"57", x"2f", x"04", x"e7",
    x"cf", x"ed", x"e4", x"d2", x"f8", x"f1", x"e3", x"d2",
    x"e0", x"e1", x"04", x"c7", x"fa", x"19", x"0d", x"fa",
    x"49", x"ed", x"ec", x"c5", x"f7", x"f5", x"12", x"06",
    x"21", x"fb", x"f8", x"16", x"23", x"00", x"d4", x"22",
    x"2f", x"ef", x"25", x"ee", x"19", x"d9", x"15", x"10",
    x"d9", x"00", x"b9", x"13", x"f7", x"18", x"fc", x"f5",
    x"15", x"92", x"d1", x"23", x"16", x"0c", x"20", x"da",
    x"35", x"05", x"cc", x"16", x"2b", x"f1", x"0d", x"f1",
    x"be", x"12", x"14", x"d8", x"d4", x"14", x"ea", x"10",
    x"3e", x"c5", x"ba", x"04", x"1f", x"d9", x"25", x"01",
    x"06", x"fd", x"fd", x"fc", x"ff", x"04", x"05", x"06",
    x"cd", x"f6", x"eb", x"96", x"2b", x"17", x"0e", x"0e",
    x"fd", x"fb", x"01", x"ff", x"fa", x"00", x"fc", x"fa",
    x"06", x"05", x"e3", x"62", x"b3", x"1b", x"e8", x"f9",
    x"13", x"03", x"d9", x"22", x"00", x"f0", x"2e", x"c8",
    x"9e", x"26", x"00", x"f9", x"06", x"3d", x"11", x"f5",
    x"0c", x"f6", x"af", x"d5", x"f0", x"07", x"b3", x"ce",
    x"20", x"29", x"0e", x"33", x"1d", x"37", x"24", x"05",
    x"f6", x"00", x"d6", x"18", x"ef", x"d3", x"0d", x"63",
    x"e1", x"e2", x"d3", x"bf", x"38", x"4d", x"dd", x"1e",
    x"40", x"42", x"2a", x"29", x"09", x"20", x"b3", x"cb",
    x"f6", x"1b", x"1e", x"e7", x"17", x"07", x"ef", x"e3",
    x"09", x"08", x"f8", x"da", x"22", x"d9", x"d2", x"26",
    x"24", x"dc", x"29", x"97", x"f5", x"0a", x"f1", x"00",
    x"12", x"de", x"f3", x"2a", x"e9", x"18", x"08", x"cf",
    x"d2", x"ff", x"00", x"b6", x"5e", x"f0", x"c9", x"11",
    x"1f", x"c2", x"fd", x"e4", x"45", x"f4", x"4d", x"fd",
    x"a1", x"52", x"df", x"d5", x"00", x"28", x"f1", x"e2",
    x"91", x"0a", x"0b", x"05", x"f8", x"f1", x"03", x"0b",
    x"22", x"d4", x"fa", x"05", x"2b", x"e7", x"f6", x"06",
    x"d9", x"19", x"f7", x"1f", x"00", x"cf", x"f8", x"f2",
    x"0c", x"23", x"15", x"bf", x"ad", x"38", x"19", x"f4",
    x"fa", x"2c", x"ea", x"b5", x"e0", x"44", x"b0", x"0b",
    x"24", x"05", x"d7", x"f1", x"f2", x"e6", x"d0", x"34",
    x"17", x"00", x"4f", x"fa", x"32", x"3f", x"e9", x"f7",
    x"f5", x"e3", x"fa", x"29", x"1d", x"d5", x"ee", x"d8",
    x"fd", x"e4", x"dd", x"ae", x"01", x"12", x"dd", x"0c",
    x"da", x"f4", x"c0", x"e9", x"20", x"2b", x"15", x"18",
    x"e3", x"13", x"3a", x"0f", x"ed", x"09", x"36", x"0e",
    x"e9", x"59", x"fa", x"ef", x"4a", x"41", x"f2", x"49",
    x"f6", x"02", x"e6", x"f4", x"e2", x"40", x"ea", x"de",
    x"ed", x"19", x"7a", x"e1", x"fc", x"0b", x"3c", x"92",
    x"e0", x"53", x"34", x"f3", x"ef", x"09", x"27", x"ae",
    x"db", x"13", x"1f", x"0d", x"ff", x"b6", x"ef", x"1b",
    x"d2", x"ce", x"06", x"ad", x"f1", x"34", x"84", x"db",
    x"ef", x"29", x"15", x"e2", x"6e", x"35", x"50", x"fe",
    x"07", x"fe", x"02", x"f9", x"fe", x"02", x"03", x"02",
    x"d9", x"fa", x"fd", x"5c", x"0e", x"f8", x"fe", x"eb",
    x"dc", x"05", x"fb", x"fc", x"fa", x"05", x"02", x"07",
    x"01", x"07", x"e8", x"03", x"12", x"41", x"2c", x"13",
    x"c8", x"1e", x"f8", x"d9", x"c4", x"e4", x"0a", x"13",
    x"1a", x"e2", x"eb", x"97", x"e1", x"d2", x"0c", x"bd",
    x"6a", x"d9", x"56", x"c7", x"f7", x"84", x"1d", x"25",
    x"f0", x"e6", x"21", x"06", x"f1", x"21", x"c4", x"e2",
    x"03", x"d7", x"1f", x"f6", x"3c", x"f7", x"0a", x"07",
    x"2d", x"08", x"a0", x"de", x"f5", x"17", x"f6", x"4b",
    x"0d", x"0b", x"10", x"88", x"f1", x"9a", x"0c", x"3a",
    x"23", x"c2", x"e2", x"0b", x"e6", x"e3", x"26", x"b3",
    x"d3", x"26", x"e9", x"be", x"37", x"ba", x"da", x"f9",
    x"04", x"1e", x"35", x"a1", x"0b", x"1a", x"01", x"27",
    x"ed", x"25", x"12", x"13", x"3d", x"30", x"fe", x"f2",
    x"a5", x"f1", x"10", x"f7", x"0c", x"26", x"d4", x"d8",
    x"09", x"e5", x"31", x"62", x"1d", x"27", x"8a", x"b5",
    x"2a", x"d7", x"1c", x"ce", x"11", x"d2", x"df", x"f5",
    x"2b", x"2c", x"0c", x"e7", x"1a", x"07", x"05", x"fd",
    x"63", x"03", x"f0", x"08", x"ce", x"d4", x"2c", x"1b",
    x"37", x"d3", x"e9", x"f8", x"10", x"f0", x"c2", x"3b",
    x"eb", x"d8", x"19", x"25", x"10", x"e0", x"fa", x"0d",
    x"15", x"a0", x"0f", x"ce", x"f7", x"28", x"e4", x"df",
    x"fb", x"11", x"f9", x"20", x"a9", x"45", x"49", x"d1",
    x"be", x"e8", x"dc", x"b3", x"29", x"e4", x"1f", x"f7",
    x"ff", x"07", x"25", x"fa", x"1e", x"1d", x"fd", x"d0",
    x"d9", x"f8", x"c6", x"ba", x"e6", x"d6", x"fd", x"fe",
    x"0c", x"17", x"aa", x"0d", x"17", x"f9", x"30", x"44",
    x"df", x"b2", x"c2", x"c3", x"1e", x"c6", x"24", x"09",
    x"b5", x"b6", x"1a", x"a2", x"f8", x"b7", x"86", x"09",
    x"f5", x"e6", x"e8", x"5f", x"66", x"ee", x"00", x"ff",
    x"ed", x"8f", x"f0", x"ef", x"a4", x"25", x"e6", x"cb",
    x"95", x"af", x"d6", x"fa", x"fd", x"b5", x"82", x"f2",
    x"c6", x"be", x"07", x"11", x"ea", x"c7", x"aa", x"21",
    x"05", x"d9", x"95", x"e7", x"cc", x"b4", x"04", x"bd",
    x"c3", x"1c", x"0f", x"ee", x"04", x"1b", x"e9", x"06",
    x"01", x"fc", x"f9", x"01", x"fa", x"01", x"06", x"fb",
    x"55", x"0a", x"e6", x"19", x"0f", x"a8", x"27", x"56",
    x"35", x"03", x"05", x"00", x"03", x"05", x"07", x"fc",
    x"05", x"fb", x"c3", x"f4", x"5c", x"b9", x"e9", x"f2",
    x"06", x"ba", x"b1", x"15", x"53", x"b8", x"f4", x"24",
    x"74", x"18", x"13", x"1d", x"e1", x"c5", x"c6", x"e5",
    x"82", x"b4", x"df", x"ae", x"9f", x"19", x"6c", x"bd",
    x"00", x"e5", x"8d", x"02", x"f7", x"09", x"11", x"20",
    x"0e", x"0b", x"ec", x"0f", x"ea", x"dc", x"ce", x"67",
    x"6e", x"ef", x"d6", x"10", x"d4", x"c9", x"b2", x"84",
    x"5a", x"e0", x"b1", x"07", x"d4", x"d3", x"f7", x"e9",
    x"27", x"e5", x"cb", x"b2", x"0c", x"cc", x"d2", x"18",
    x"f1", x"a5", x"85", x"a4", x"12", x"cd", x"78", x"68",
    x"0f", x"fe", x"8a", x"2b", x"33", x"f7", x"15", x"2d",
    x"20", x"fb", x"2f", x"fe", x"01", x"00", x"c8", x"26",
    x"f7", x"c1", x"32", x"f8", x"13", x"22", x"ff", x"05",
    x"1f", x"08", x"e5", x"1b", x"31", x"0d", x"fc", x"f1",
    x"bf", x"0d", x"04", x"ff", x"ec", x"f0", x"eb", x"18",
    x"22", x"13", x"38", x"07", x"08", x"30", x"60", x"68",
    x"f5", x"cd", x"b4", x"9d", x"60", x"aa", x"b7", x"b9",
    x"fd", x"15", x"c9", x"b0", x"2c", x"f0", x"f6", x"1d",
    x"22", x"10", x"eb", x"f0", x"e6", x"f1", x"17", x"da",
    x"0f", x"00", x"85", x"03", x"14", x"9d", x"fe", x"cb",
    x"72", x"2d", x"e7", x"b1", x"ed", x"e8", x"16", x"15",
    x"fa", x"e1", x"e0", x"f8", x"e2", x"a7", x"20", x"a2",
    x"b2", x"fb", x"34", x"f8", x"f0", x"8b", x"fd", x"0e",
    x"0b", x"ca", x"ed", x"f7", x"d3", x"c7", x"e5", x"7c",
    x"f9", x"17", x"ec", x"9c", x"97", x"0e", x"d3", x"a3",
    x"ee", x"5d", x"39", x"d9", x"05", x"41", x"a8", x"98",
    x"83", x"08", x"14", x"e1", x"bb", x"0e", x"0a", x"ff",
    x"11", x"c0", x"1a", x"21", x"2e", x"2e", x"16", x"28",
    x"fd", x"08", x"17", x"2f", x"0a", x"62", x"ea", x"e0",
    x"c5", x"d3", x"c2", x"b0", x"23", x"0f", x"9e", x"10",
    x"2c", x"1e", x"f0", x"23", x"1a", x"4a", x"dc", x"f3",
    x"e7", x"b5", x"d0", x"c7", x"b9", x"d6", x"c1", x"de",
    x"e6", x"d7", x"01", x"ce", x"36", x"0a", x"02", x"fa",
    x"03", x"04", x"05", x"f9", x"fe", x"00", x"03", x"fb",
    x"d9", x"dc", x"24", x"00", x"12", x"f9", x"14", x"0b",
    x"af", x"fc", x"fa", x"04", x"07", x"05", x"fd", x"fd",
    x"02", x"02", x"d5", x"cc", x"bc", x"0b", x"ef", x"43",
    x"3d", x"07", x"4c", x"10", x"1c", x"64", x"f4", x"f8",
    x"cc", x"e6", x"11", x"fd", x"a4", x"f8", x"dc", x"ce",
    x"32", x"e7", x"18", x"f1", x"f9", x"36", x"0e", x"ee",
    x"24", x"17", x"03", x"23", x"47", x"f8", x"17", x"ef",
    x"f5", x"14", x"fd", x"1f", x"00", x"cd", x"f5", x"02",
    x"d1", x"c4", x"d1", x"08", x"f8", x"e8", x"ec", x"ee",
    x"f8", x"f7", x"00", x"20", x"d0", x"22", x"1d", x"0d",
    x"24", x"18", x"ec", x"e1", x"04", x"fe", x"24", x"4b",
    x"d8", x"37", x"23", x"11", x"49", x"d3", x"c2", x"60",
    x"36", x"03", x"f2", x"ec", x"04", x"fb", x"91", x"ee",
    x"fb", x"b8", x"0c", x"36", x"53", x"f5", x"19", x"f5",
    x"05", x"ec", x"f3", x"08", x"0c", x"09", x"09", x"e7",
    x"f4", x"46", x"2f", x"1a", x"35", x"0e", x"a8", x"1a",
    x"0b", x"90", x"02", x"1f", x"e6", x"3a", x"06", x"f5",
    x"15", x"0e", x"fb", x"01", x"37", x"06", x"e1", x"0f",
    x"fa", x"14", x"ec", x"30", x"fb", x"e3", x"29", x"17",
    x"cd", x"b8", x"ca", x"c9", x"b9", x"08", x"00", x"fe",
    x"09", x"07", x"fc", x"ca", x"db", x"21", x"1a", x"31",
    x"16", x"f7", x"f7", x"2d", x"2c", x"48", x"52", x"be",
    x"4e", x"bc", x"d2", x"fd", x"dc", x"0c", x"94", x"c6",
    x"2d", x"26", x"02", x"0e", x"d0", x"4b", x"27", x"40",
    x"06", x"1a", x"3d", x"f8", x"ec", x"8a", x"ed", x"f1",
    x"fb", x"e2", x"d9", x"e4", x"db", x"09", x"d6", x"28",
    x"f2", x"b4", x"0c", x"c7", x"d7", x"0b", x"26", x"3c",
    x"24", x"01", x"ee", x"0e", x"12", x"1d", x"e7", x"25",
    x"19", x"ed", x"d8", x"d6", x"ea", x"e8", x"eb", x"de",
    x"01", x"26", x"03", x"d9", x"ed", x"df", x"fc", x"18",
    x"a8", x"e6", x"9e", x"1f", x"20", x"2f", x"38", x"06",
    x"4c", x"00", x"36", x"58", x"17", x"46", x"0b", x"10",
    x"d2", x"08", x"23", x"a6", x"67", x"e2", x"e5", x"15",
    x"1f", x"fc", x"f8", x"ed", x"25", x"e9", x"03", x"e5",
    x"e8", x"d7", x"f8", x"13", x"f5", x"f8", x"0c", x"f9",
    x"fa", x"ff", x"ff", x"fb", x"05", x"06", x"fa", x"06",
    x"06", x"18", x"2a", x"27", x"d1", x"e5", x"22", x"62",
    x"39", x"fa", x"fc", x"fa", x"01", x"04", x"02", x"00",
    x"fd", x"02", x"2a", x"0a", x"a8", x"25", x"27", x"0d",
    x"32", x"f8", x"e7", x"4b", x"cd", x"04", x"01", x"3d",
    x"f2", x"12", x"0e", x"ae", x"17", x"df", x"0c", x"35",
    x"e6", x"f3", x"dd", x"09", x"e7", x"f1", x"fc", x"18",
    x"51", x"4f", x"38", x"22", x"fd", x"e1", x"11", x"fc",
    x"fa", x"39", x"0b", x"b3", x"26", x"3b", x"e6", x"9c",
    x"02", x"20", x"5d", x"02", x"fb", x"e0", x"52", x"2f",
    x"eb", x"cd", x"0d", x"f1", x"fa", x"19", x"e9", x"17",
    x"f6", x"1c", x"de", x"8b", x"03", x"ac", x"dd", x"19",
    x"d5", x"70", x"30", x"dd", x"ef", x"48", x"21", x"1c",
    x"f6", x"37", x"15", x"e2", x"0a", x"22", x"f4", x"09",
    x"e5", x"64", x"2c", x"d2", x"cf", x"d4", x"4c", x"14",
    x"17", x"07", x"05", x"13", x"ec", x"1c", x"db", x"e4",
    x"f9", x"dc", x"0a", x"16", x"fd", x"f5", x"e0", x"fd",
    x"06", x"47", x"10", x"d6", x"fa", x"e3", x"d9", x"f9",
    x"f0", x"53", x"fb", x"d1", x"ff", x"ee", x"d7", x"46",
    x"f5", x"db", x"d4", x"47", x"0d", x"5c", x"08", x"38",
    x"3f", x"14", x"e9", x"07", x"00", x"00", x"f6", x"1a",
    x"33", x"fc", x"ec", x"e2", x"e5", x"08", x"dd", x"08",
    x"14", x"c6", x"8f", x"03", x"27", x"2a", x"1a", x"11",
    x"df", x"14", x"f0", x"21", x"de", x"1f", x"13", x"40",
    x"da", x"df", x"df", x"e6", x"dd", x"28", x"f2", x"fc",
    x"03", x"f1", x"47", x"03", x"32", x"42", x"e4", x"a9",
    x"d4", x"9e", x"ff", x"ed", x"b9", x"a2", x"f4", x"ec",
    x"32", x"1f", x"11", x"eb", x"0d", x"d3", x"ea", x"29",
    x"0d", x"19", x"33", x"d1", x"0c", x"40", x"ea", x"dd",
    x"12", x"06", x"04", x"21", x"2a", x"f5", x"1d", x"89",
    x"20", x"23", x"06", x"1d", x"0f", x"e7", x"32", x"4f",
    x"08", x"22", x"07", x"fe", x"1f", x"0e", x"fb", x"11",
    x"f2", x"10", x"1c", x"0a", x"d3", x"e1", x"d8", x"12",
    x"ed", x"fc", x"cb", x"c1", x"c0", x"05", x"19", x"ff",
    x"cb", x"14", x"35", x"bf", x"e3", x"e9", x"fc", x"fd",
    x"19", x"db", x"13", x"17", x"2d", x"f9", x"2a", x"f9",
    x"00", x"07", x"fe", x"07", x"06", x"02", x"06", x"fa",
    x"cf", x"dd", x"d5", x"d9", x"a0", x"ec", x"d7", x"21",
    x"ed", x"03", x"fb", x"fb", x"ff", x"fa", x"01", x"01",
    x"ff", x"01", x"d2", x"e6", x"0a", x"d0", x"bb", x"24",
    x"16", x"15", x"0b", x"df", x"d1", x"29", x"e7", x"cb",
    x"19", x"3f", x"09", x"03", x"00", x"2a", x"14", x"ed",
    x"3c", x"08", x"db", x"e4", x"d4", x"ff", x"f9", x"fa",
    x"de", x"d8", x"ea", x"df", x"5d", x"f5", x"ef", x"c9",
    x"f8", x"47", x"e5", x"e3", x"fb", x"e3", x"c1", x"6a",
    x"3b", x"15", x"ea", x"21", x"0f", x"b8", x"06", x"bb",
    x"08", x"43", x"21", x"09", x"3b", x"49", x"fe", x"fe",
    x"2f", x"ff", x"0c", x"0e", x"ff", x"03", x"0a", x"13",
    x"fa", x"db", x"08", x"37", x"1b", x"db", x"15", x"08",
    x"f5", x"1c", x"ee", x"b7", x"0d", x"16", x"4f", x"ed",
    x"12", x"16", x"f2", x"1b", x"10", x"17", x"0d", x"da",
    x"17", x"01", x"f9", x"eb", x"0d", x"e3", x"20", x"21",
    x"01", x"eb", x"f7", x"02", x"df", x"f9", x"f8", x"fa",
    x"0a", x"9b", x"9d", x"e9", x"76", x"c2", x"af", x"02",
    x"f6", x"bb", x"dd", x"ec", x"bb", x"bb", x"f8", x"1b",
    x"f8", x"ea", x"1e", x"e8", x"d7", x"e1", x"82", x"14",
    x"0f", x"db", x"f0", x"32", x"f1", x"d9", x"1b", x"e4",
    x"fa", x"e1", x"e1", x"d3", x"0a", x"16", x"e1", x"05",
    x"d7", x"03", x"24", x"c7", x"ff", x"10", x"d8", x"f7",
    x"3b", x"ec", x"fa", x"10", x"0a", x"14", x"0e", x"c2",
    x"b4", x"22", x"55", x"83", x"b6", x"eb", x"26", x"26",
    x"fa", x"2d", x"1c", x"e9", x"1f", x"1f", x"05", x"e1",
    x"16", x"06", x"ce", x"0a", x"09", x"e3", x"05", x"03",
    x"24", x"f7", x"fd", x"54", x"06", x"f0", x"fb", x"e7",
    x"15", x"09", x"e1", x"2b", x"fd", x"17", x"13", x"b3",
    x"f1", x"07", x"00", x"49", x"2b", x"2d", x"19", x"e6",
    x"e6", x"11", x"f1", x"cd", x"f0", x"c8", x"f7", x"2b",
    x"2f", x"21", x"14", x"39", x"09", x"2a", x"1d", x"fd",
    x"3d", x"29", x"6b", x"2b", x"e9", x"e8", x"0d", x"00",
    x"23", x"41", x"c8", x"00", x"e9", x"12", x"01", x"ff",
    x"e2", x"d5", x"05", x"31", x"1c", x"13", x"0f", x"dd",
    x"c8", x"37", x"ef", x"fe", x"9b", x"18", x"05", x"01",
    x"f9", x"fc", x"03", x"02", x"04", x"fd", x"07", x"f9",
    x"2a", x"2c", x"40", x"f3", x"bb", x"bc", x"cc", x"e6",
    x"c8", x"f9", x"01", x"fa", x"fd", x"02", x"02", x"ff",
    x"fe", x"fb", x"fb", x"05", x"1d", x"f8", x"1b", x"19",
    x"f0", x"1f", x"27", x"c9", x"15", x"f5", x"35", x"24",
    x"3c", x"59", x"1e", x"10", x"43", x"e1", x"ed", x"2a",
    x"0d", x"ef", x"e3", x"31", x"0e", x"33", x"1f", x"0c",
    x"24", x"c3", x"e5", x"e1", x"3c", x"43", x"0a", x"16",
    x"e1", x"e8", x"ed", x"40", x"c1", x"4c", x"3d", x"19",
    x"fc", x"df", x"1b", x"0f", x"18", x"0b", x"25", x"45",
    x"26", x"e5", x"05", x"07", x"f7", x"e0", x"f3", x"46",
    x"e6", x"30", x"0e", x"3c", x"d7", x"e7", x"07", x"09",
    x"14", x"21", x"f5", x"d2", x"13", x"17", x"e6", x"17",
    x"e8", x"00", x"fb", x"d5", x"06", x"fd", x"21", x"20",
    x"41", x"8c", x"c7", x"93", x"cf", x"ca", x"16", x"fb",
    x"af", x"ce", x"12", x"a8", x"b1", x"33", x"1b", x"0f",
    x"fb", x"ec", x"03", x"4a", x"e4", x"22", x"20", x"15",
    x"f9", x"35", x"08", x"f5", x"1d", x"be", x"f4", x"e1",
    x"19", x"de", x"d7", x"b8", x"1e", x"f7", x"08", x"34",
    x"28", x"26", x"0c", x"01", x"fe", x"df", x"ef", x"85",
    x"3c", x"05", x"ec", x"de", x"58", x"17", x"e4", x"70",
    x"88", x"03", x"1b", x"e6", x"fb", x"ec", x"f9", x"08",
    x"0d", x"2d", x"46", x"f6", x"db", x"f7", x"2a", x"fe",
    x"4e", x"dc", x"e4", x"21", x"04", x"ee", x"07", x"0f",
    x"23", x"05", x"21", x"35", x"f2", x"f5", x"fb", x"0a",
    x"3d", x"0d", x"0f", x"0c", x"dc", x"e6", x"f1", x"b5",
    x"c7", x"cb", x"d0", x"76", x"e7", x"ec", x"03", x"ff",
    x"ca", x"de", x"12", x"f2", x"2e", x"f0", x"0d", x"0e",
    x"e3", x"e3", x"01", x"bd", x"e6", x"b9", x"91", x"9e",
    x"c6", x"2c", x"f1", x"1a", x"4a", x"e0", x"f5", x"03",
    x"0c", x"c7", x"d9", x"d0", x"0a", x"2a", x"ec", x"2b",
    x"12", x"2d", x"4a", x"d6", x"f3", x"f4", x"c6", x"e0",
    x"ba", x"0c", x"09", x"f8", x"39", x"ed", x"22", x"23",
    x"0e", x"fa", x"26", x"03", x"fb", x"e2", x"77", x"09",
    x"db", x"c2", x"17", x"0b", x"18", x"28", x"dd", x"b1",
    x"a1", x"12", x"1b", x"e7", x"1f", x"22", x"08", x"f9",
    x"fd", x"05", x"01", x"f9", x"05", x"01", x"00", x"fa",
    x"ce", x"e3", x"32", x"ff", x"07", x"16", x"f6", x"fa",
    x"e9", x"07", x"05", x"fb", x"fc", x"04", x"07", x"fa",
    x"f9", x"fd", x"fe", x"29", x"0c", x"fd", x"54", x"2b",
    x"f1", x"21", x"29", x"ef", x"f8", x"dd", x"f6", x"0c",
    x"32", x"19", x"c1", x"ed", x"e2", x"e4", x"d5", x"e3",
    x"02", x"f5", x"3f", x"28", x"04", x"27", x"08", x"28",
    x"04", x"ec", x"fb", x"01", x"f5", x"06", x"df", x"3e",
    x"00", x"f3", x"0b", x"c9", x"05", x"f0", x"2e", x"35",
    x"f2", x"bc", x"26", x"ff", x"07", x"34", x"fd", x"1c",
    x"9b", x"0e", x"0f", x"f6", x"f6", x"d0", x"d7", x"36",
    x"3d", x"f4", x"a9", x"eb", x"2e", x"f7", x"29", x"31",
    x"f8", x"62", x"a3", x"7e", x"c1", x"c1", x"d7", x"77",
    x"2b", x"ee", x"00", x"38", x"ff", x"f6", x"10", x"1c",
    x"1e", x"30", x"21", x"08", x"05", x"9b", x"3a", x"3e",
    x"d5", x"cb", x"0e", x"2e", x"01", x"24", x"12", x"09",
    x"14", x"28", x"24", x"24", x"01", x"00", x"eb", x"ec",
    x"19", x"11", x"3b", x"40", x"3a", x"fa", x"df", x"f3",
    x"68", x"2b", x"0c", x"15", x"46", x"22", x"f1", x"32",
    x"31", x"f0", x"2d", x"1b", x"bc", x"03", x"22", x"ca",
    x"44", x"ca", x"87", x"be", x"ff", x"ea", x"00", x"02",
    x"b9", x"bb", x"db", x"49", x"56", x"0a", x"08", x"4b",
    x"3e", x"ba", x"20", x"27", x"0b", x"ec", x"f2", x"d4",
    x"d9", x"bc", x"e8", x"17", x"ec", x"e3", x"21", x"fe",
    x"f4", x"f9", x"28", x"eb", x"ed", x"f3", x"f1", x"69",
    x"fd", x"14", x"32", x"bb", x"fe", x"f7", x"f4", x"ef",
    x"d6", x"e5", x"b8", x"ff", x"e8", x"cf", x"dd", x"1a",
    x"13", x"b5", x"1b", x"bc", x"af", x"f3", x"f0", x"12",
    x"37", x"d1", x"48", x"d9", x"2a", x"2f", x"fc", x"0d",
    x"36", x"a0", x"ac", x"25", x"c2", x"fb", x"31", x"ff",
    x"06", x"31", x"f7", x"f1", x"3a", x"0a", x"38", x"ee",
    x"1c", x"18", x"89", x"d2", x"4f", x"f0", x"36", x"03",
    x"36", x"13", x"1c", x"df", x"c5", x"70", x"62", x"0c",
    x"f4", x"0a", x"f3", x"c7", x"bc", x"5b", x"ca", x"0e",
    x"17", x"16", x"14", x"05", x"c4", x"58", x"04", x"fa",
    x"14", x"00", x"1d", x"e2", x"1d", x"eb", x"f4", x"fc",
    x"06", x"05", x"fa", x"00", x"03", x"05", x"06", x"04",
    x"17", x"f9", x"11", x"eb", x"e2", x"f8", x"2c", x"f6",
    x"12", x"06", x"fd", x"fb", x"01", x"f9", x"fd", x"ff",
    x"06", x"f9", x"e6", x"91", x"2c", x"bb", x"0f", x"2c",
    x"25", x"28", x"21", x"d4", x"cb", x"17", x"96", x"df",
    x"db", x"f1", x"fe", x"f8", x"c6", x"fa", x"2b", x"f9",
    x"0b", x"0b", x"0e", x"0b", x"11", x"16", x"00", x"58",
    x"07", x"f8", x"1f", x"46", x"20", x"c5", x"4b", x"90",
    x"e1", x"bf", x"f0", x"ad", x"fe", x"1b", x"ea", x"57",
    x"73", x"89", x"32", x"fa", x"25", x"21", x"01", x"f1",
    x"12", x"27", x"66", x"1c", x"38", x"0d", x"f0", x"a7",
    x"9f", x"39", x"12", x"0d", x"14", x"1a", x"04", x"1d",
    x"ae", x"48", x"f8", x"b5", x"2a", x"cd", x"36", x"5c",
    x"db", x"03", x"04", x"8b", x"1b", x"22", x"30", x"2d",
    x"11", x"f6", x"03", x"c8", x"29", x"02", x"34", x"16",
    x"35", x"3c", x"fa", x"2a", x"0b", x"fd", x"fc", x"fb",
    x"f6", x"16", x"03", x"25", x"15", x"1c", x"a0", x"20",
    x"ba", x"df", x"b9", x"f6", x"3b", x"18", x"e1", x"6d",
    x"ed", x"a0", x"23", x"5b", x"e0", x"34", x"2a", x"1a",
    x"2e", x"bf", x"c1", x"17", x"32", x"18", x"08", x"fa",
    x"f1", x"e8", x"f2", x"c8", x"e7", x"f2", x"f1", x"fc",
    x"33", x"2f", x"17", x"b3", x"de", x"fa", x"e2", x"e2",
    x"2e", x"e3", x"6c", x"ea", x"bc", x"d6", x"28", x"4b",
    x"4c", x"2f", x"03", x"14", x"64", x"c8", x"ab", x"fd",
    x"f1", x"01", x"3a", x"f6", x"dd", x"b7", x"8d", x"cd",
    x"c6", x"f7", x"35", x"e4", x"fb", x"fa", x"0f", x"ff",
    x"ec", x"be", x"d5", x"b9", x"ca", x"e2", x"d3", x"dc",
    x"c2", x"2b", x"33", x"27", x"fa", x"27", x"0f", x"1b",
    x"04", x"05", x"03", x"f6", x"03", x"fa", x"fc", x"01",
    x"ff", x"03", x"f7", x"f9", x"01", x"fb", x"fb", x"ff",
    x"f7", x"ff", x"fe", x"fe", x"fb", x"f9", x"02", x"f8",
    x"fd", x"fb", x"02", x"01", x"ff", x"fd", x"f8", x"fb",
    x"02", x"fc", x"fc", x"ff", x"fd", x"02", x"fc", x"f9",
    x"fa", x"fa", x"fd", x"f9", x"fb", x"fb", x"fa", x"03",
    x"01", x"02", x"01", x"ff", x"fc", x"04", x"01", x"fb",
    x"02", x"fa", x"00", x"f8", x"01", x"fc", x"00", x"fc",
    x"01", x"06", x"fb", x"02", x"f9", x"fb", x"fa", x"fc",
    x"f8", x"ff", x"fd", x"f9", x"02", x"f9", x"f4", x"fa",
    x"01", x"ff", x"03", x"03", x"04", x"06", x"fc", x"fb",
    x"04", x"03", x"00", x"02", x"00", x"fc", x"00", x"f9",
    x"f9", x"f7", x"fa", x"01", x"01", x"fb", x"fc", x"fc",
    x"fe", x"fa", x"fa", x"04", x"fd", x"05", x"fe", x"00",
    x"fd", x"01", x"fb", x"03", x"00", x"f5", x"f9", x"f8",
    x"f8", x"02", x"fd", x"01", x"01", x"f8", x"fb", x"01",
    x"fe", x"03", x"fc", x"fa", x"fe", x"f7", x"f6", x"fb",
    x"f8", x"fe", x"f7", x"05", x"03", x"fd", x"f7", x"04",
    x"fd", x"f9", x"01", x"04", x"04", x"fd", x"fb", x"f6",
    x"fe", x"fc", x"05", x"ff", x"ff", x"03", x"fe", x"02",
    x"fc", x"fe", x"fd", x"f9", x"f9", x"00", x"ff", x"02",
    x"fa", x"f9", x"03", x"fe", x"03", x"f9", x"00", x"01",
    x"01", x"f8", x"fa", x"01", x"01", x"06", x"fd", x"01",
    x"00", x"fe", x"fd", x"fe", x"f9", x"02", x"fa", x"02",
    x"f9", x"02", x"fb", x"fa", x"fc", x"f6", x"ff", x"fe",
    x"05", x"ff", x"fe", x"ff", x"fd", x"fa", x"fc", x"fb",
    x"f8", x"04", x"fa", x"f9", x"05", x"f9", x"f6", x"02",
    x"fa", x"f9", x"02", x"fb", x"f8", x"f9", x"ff", x"fe",
    x"05", x"f9", x"01", x"02", x"f5", x"05", x"ff", x"f7",
    x"02", x"f6", x"f9", x"fc", x"f6", x"fa", x"01", x"ff",
    x"f8", x"f8", x"f4", x"04", x"01", x"f7", x"ff", x"05",
    x"fb", x"fd", x"01", x"04", x"fe", x"03", x"fd", x"f8",
    x"f5", x"fd", x"f8", x"fb", x"00", x"03", x"f8", x"05",
    x"fe", x"fd", x"ff", x"ff", x"fc", x"fb", x"03", x"fb",
    x"f6", x"f5", x"f6", x"fe", x"fd", x"01", x"f8", x"fb",
    x"f7", x"fb", x"f5", x"f3", x"f5", x"fe", x"02", x"f5",
    x"22", x"20", x"1d", x"1a", x"17", x"13", x"a9", x"ad",
    x"9f", x"35", x"19", x"2e", x"2c", x"fd", x"f6", x"ee",
    x"e7", x"f6", x"bc", x"d0", x"f8", x"07", x"1a", x"ff",
    x"e2", x"ba", x"4a", x"29", x"e6", x"21", x"c2", x"1a",
    x"36", x"e7", x"33", x"3d", x"3c", x"03", x"0e", x"13",
    x"25", x"2e", x"a6", x"df", x"b0", x"f7", x"d7", x"1b",
    x"d6", x"ea", x"10", x"00", x"d4", x"c0", x"e3", x"fa",
    x"e7", x"cf", x"0e", x"76", x"94", x"98", x"7f", x"f9",
    x"fc", x"fc", x"fc", x"f9", x"f9", x"fb", x"03", x"02",
    x"59", x"e2", x"f1", x"da", x"8d", x"a6", x"29", x"02",
    x"a1", x"fa", x"01", x"04", x"07", x"00", x"ff", x"01",
    x"02", x"fa", x"17", x"14", x"ed", x"32", x"0b", x"ea",
    x"a6", x"db", x"de", x"ec", x"f5", x"00", x"4d", x"21",
    x"21", x"74", x"b3", x"fe", x"18", x"01", x"09", x"c4",
    x"fb", x"f5", x"b5", x"1e", x"29", x"11", x"15", x"12",
    x"d5", x"06", x"41", x"be", x"26", x"2b", x"ee", x"f5",
    x"08", x"74", x"2d", x"14", x"db", x"fb", x"99", x"fd",
    x"ff", x"3d", x"dc", x"03", x"08", x"c7", x"48", x"3a",
    x"e5", x"d4", x"eb", x"b8", x"b0", x"8f", x"e9", x"be",
    x"7c", x"ff", x"eb", x"ee", x"09", x"ec", x"db", x"18",
    x"fa", x"c7", x"28", x"0e", x"2b", x"fe", x"f4", x"f6",
    x"f5", x"f6", x"ca", x"07", x"4b", x"fa", x"02", x"dd",
    x"c2", x"f7", x"5d", x"52", x"3b", x"15", x"19", x"a9",
    x"a4", x"05", x"e0", x"49", x"c0", x"45", x"02", x"1b",
    x"f1", x"a1", x"04", x"8c", x"eb", x"0a", x"2d", x"ec",
    x"15", x"a2", x"70", x"eb", x"3e", x"e9", x"da", x"0c",
    x"e5", x"07", x"d4", x"09", x"fb", x"0a", x"d5", x"fc",
    x"ff", x"20", x"07", x"36", x"1e", x"e2", x"04", x"1a",
    x"d8", x"29", x"f9", x"f4", x"0e", x"fe", x"bc", x"76",
    x"d8", x"17", x"1c", x"fc", x"1e", x"0c", x"fc", x"f7",
    x"f3", x"03", x"d2", x"44", x"20", x"39", x"03", x"09",
    x"08", x"9d", x"c1", x"79", x"2d", x"26", x"27", x"ae",
    x"f2", x"15", x"06", x"32", x"00", x"0e", x"00", x"0e",
    x"33", x"0a", x"11", x"cf", x"d7", x"f6", x"f7", x"cb",
    x"d9", x"04", x"f2", x"ee", x"fb", x"0c", x"f4", x"0f",
    x"11", x"33", x"f3", x"f6", x"12", x"e1", x"ee", x"2e",
    x"05", x"2d", x"dc", x"42", x"21", x"d8", x"df", x"f1",
    x"30", x"0c", x"45", x"1b", x"ca", x"15", x"1a", x"e3",
    x"fc", x"18", x"d7", x"2d", x"d6", x"e9", x"11", x"19",
    x"13", x"1d", x"14", x"22", x"20", x"e7", x"5a", x"0a",
    x"ee", x"26", x"4a", x"e8", x"a0", x"86", x"de", x"ef",
    x"0f", x"d1", x"0f", x"39", x"02", x"8f", x"7a", x"dd",
    x"d3", x"c3", x"ac", x"e9", x"0e", x"d9", x"d8", x"e6",
    x"db", x"f6", x"00", x"1e", x"d0", x"db", x"f3", x"06",
    x"05", x"ff", x"f9", x"00", x"fb", x"00", x"03", x"05",
    x"27", x"58", x"48", x"25", x"12", x"cf", x"25", x"11",
    x"fa", x"fa", x"05", x"fe", x"fe", x"fc", x"03", x"07",
    x"07", x"04", x"3a", x"1a", x"3e", x"29", x"0b", x"41",
    x"08", x"4c", x"2f", x"b9", x"e4", x"ef", x"43", x"0e",
    x"30", x"b1", x"18", x"21", x"1f", x"b3", x"84", x"10",
    x"24", x"dc", x"11", x"2f", x"14", x"be", x"f0", x"ca",
    x"f5", x"14", x"0f", x"0c", x"2a", x"17", x"37", x"ff",
    x"cf", x"23", x"16", x"e4", x"cd", x"07", x"1a", x"22",
    x"00", x"b2", x"48", x"09", x"a5", x"3d", x"35", x"c5",
    x"da", x"c1", x"cc", x"1f", x"18", x"ea", x"fa", x"03",
    x"22", x"d4", x"24", x"db", x"17", x"f8", x"e7", x"09",
    x"2b", x"15", x"2d", x"f8", x"de", x"34", x"e3", x"14",
    x"15", x"ef", x"20", x"13", x"be", x"e9", x"19", x"0b",
    x"18", x"c6", x"e7", x"c7", x"0a", x"05", x"04", x"06",
    x"04", x"14", x"04", x"0d", x"09", x"fb", x"fe", x"d4",
    x"19", x"ff", x"ea", x"03", x"f2", x"eb", x"f5", x"af",
    x"fa", x"e1", x"e6", x"d5", x"03", x"21", x"15", x"f8",
    x"f7", x"0e", x"fe", x"38", x"e0", x"c1", x"0d", x"e8",
    x"fb", x"ad", x"e8", x"18", x"17", x"f3", x"1a", x"0a",
    x"0f", x"32", x"07", x"f8", x"eb", x"30", x"2e", x"ed",
    x"f2", x"36", x"b9", x"f1", x"f6", x"dc", x"e3", x"be",
    x"04", x"1c", x"1e", x"01", x"44", x"d7", x"02", x"0b",
    x"23", x"95", x"ca", x"1e", x"c3", x"7a", x"89", x"d9",
    x"c8", x"73", x"1b", x"26", x"f9", x"09", x"ff", x"0d",
    x"26", x"e0", x"f4", x"eb", x"49", x"1d", x"ee", x"04",
    x"da", x"e2", x"df", x"03", x"f1", x"1a", x"ec", x"d7",
    x"23", x"10", x"eb", x"d7", x"f3", x"88", x"a4", x"0d",
    x"11", x"f8", x"bc", x"14", x"08", x"2f", x"00", x"04",
    x"e0", x"0b", x"fd", x"d2", x"05", x"19", x"02", x"fe",
    x"ec", x"3e", x"13", x"17", x"8c", x"76", x"e7", x"d4",
    x"fd", x"04", x"07", x"ef", x"2e", x"2e", x"eb", x"49",
    x"3c", x"a6", x"17", x"1e", x"9f", x"d3", x"cd", x"c9",
    x"e6", x"f8", x"b4", x"ce", x"f9", x"f9", x"19", x"18",
    x"0f", x"63", x"96", x"02", x"f4", x"d2", x"13", x"d2",
    x"8c", x"e4", x"e2", x"19", x"e6", x"f3", x"14", x"f9",
    x"04", x"fe", x"06", x"fa", x"04", x"fa", x"00", x"02",
    x"0f", x"33", x"c6", x"13", x"2f", x"2b", x"d2", x"1f",
    x"2c", x"06", x"01", x"00", x"ff", x"00", x"04", x"05",
    x"05", x"01", x"f1", x"4f", x"33", x"e8", x"0d", x"cb",
    x"87", x"1a", x"ec", x"9b", x"a5", x"af", x"f6", x"fa",
    x"20", x"ae", x"fa", x"f6", x"34", x"2d", x"fe", x"29",
    x"10", x"04", x"fc", x"ee", x"12", x"0b", x"1f", x"d5",
    x"dd", x"10", x"4e", x"f2", x"0f", x"2f", x"d9", x"e0",
    x"d3", x"c0", x"8f", x"1e", x"b2", x"9f", x"fc", x"3e",
    x"06", x"3b", x"0e", x"ff", x"21", x"b6", x"9c", x"00",
    x"0b", x"0f", x"a9", x"01", x"37", x"c6", x"e1", x"0f",
    x"05", x"f5", x"ed", x"fe", x"c2", x"f5", x"19", x"08",
    x"f2", x"ee", x"10", x"e8", x"cb", x"04", x"fb", x"01",
    x"f0", x"e2", x"0b", x"13", x"c9", x"25", x"13", x"bb",
    x"d0", x"d7", x"04", x"e3", x"2a", x"f5", x"13", x"d3",
    x"11", x"3d", x"fe", x"16", x"14", x"13", x"ee", x"f3",
    x"02", x"31", x"2d", x"bd", x"de", x"26", x"d4", x"f6",
    x"fd", x"e7", x"4e", x"0b", x"bf", x"8c", x"01", x"02",
    x"08", x"f2", x"a2", x"2d", x"2b", x"96", x"09", x"11",
    x"0b", x"12", x"ee", x"dc", x"23", x"0b", x"1a", x"eb",
    x"0d", x"e9", x"08", x"2a", x"f5", x"36", x"0c", x"01",
    x"fb", x"f4", x"d4", x"f4", x"c5", x"dc", x"14", x"fe",
    x"9c", x"f6", x"2b", x"fb", x"e8", x"be", x"09", x"d4",
    x"ca", x"82", x"e0", x"e9", x"ef", x"25", x"f2", x"19",
    x"12", x"12", x"d5", x"f7", x"f6", x"c3", x"d0", x"c7",
    x"fc", x"48", x"0d", x"db", x"12", x"21", x"e3", x"04",
    x"d8", x"01", x"06", x"15", x"e9", x"1f", x"1f", x"fc",
    x"c7", x"e2", x"00", x"df", x"c9", x"11", x"f4", x"2c",
    x"b8", x"cf", x"1f", x"d1", x"0a", x"e0", x"f2", x"0c",
    x"f6", x"c3", x"f8", x"fe", x"ed", x"ed", x"36", x"17",
    x"1d", x"1f", x"24", x"0e", x"fc", x"06", x"05", x"ff",
    x"cd", x"c1", x"d6", x"2b", x"fb", x"db", x"3d", x"07",
    x"03", x"1f", x"46", x"44", x"d7", x"c2", x"9d", x"34",
    x"0b", x"1e", x"18", x"01", x"06", x"f9", x"b1", x"ca",
    x"1c", x"e7", x"02", x"d9", x"02", x"fb", x"e3", x"14",
    x"09", x"f9", x"e8", x"02", x"e0", x"05", x"b3", x"fb",
    x"fe", x"fc", x"fa", x"02", x"02", x"03", x"06", x"01",
    x"66", x"1b", x"12", x"e2", x"13", x"06", x"fc", x"45",
    x"f7", x"04", x"f9", x"fe", x"05", x"fa", x"04", x"04",
    x"00", x"ff", x"2d", x"29", x"18", x"01", x"11", x"d2",
    x"2e", x"10", x"0d", x"ca", x"d1", x"d6", x"e0", x"0c",
    x"08", x"f5", x"08", x"09", x"e0", x"b9", x"b9", x"2f",
    x"08", x"34", x"32", x"4f", x"1b", x"e9", x"9c", x"04",
    x"d4", x"fc", x"1f", x"2d", x"38", x"3e", x"e4", x"c2",
    x"fc", x"0b", x"12", x"2c", x"58", x"2e", x"3b", x"1b",
    x"24", x"e9", x"17", x"e6", x"96", x"35", x"37", x"fd",
    x"fa", x"ef", x"fa", x"24", x"14", x"26", x"01", x"fa",
    x"63", x"20", x"01", x"ec", x"1b", x"f5", x"fe", x"d6",
    x"23", x"f8", x"d7", x"3e", x"63", x"28", x"0d", x"9b",
    x"fc", x"13", x"d4", x"b2", x"fe", x"e0", x"1e", x"19",
    x"ee", x"10", x"1c", x"e6", x"2a", x"04", x"03", x"e6",
    x"ee", x"ea", x"10", x"1c", x"61", x"ab", x"ec", x"0c",
    x"37", x"17", x"13", x"0e", x"ec", x"d1", x"07", x"26",
    x"09", x"d5", x"b6", x"ff", x"44", x"22", x"ef", x"f2",
    x"f9", x"c5", x"30", x"27", x"e5", x"08", x"fc", x"d8",
    x"e5", x"0b", x"f8", x"43", x"37", x"fa", x"06", x"29",
    x"03", x"8a", x"0a", x"0d", x"fb", x"17", x"42", x"e7",
    x"e8", x"f0", x"f3", x"c1", x"ee", x"f9", x"e1", x"02",
    x"20", x"25", x"35", x"b6", x"c3", x"5d", x"1d", x"0f",
    x"27", x"30", x"02", x"33", x"0a", x"c8", x"f7", x"14",
    x"01", x"15", x"19", x"0c", x"bc", x"19", x"33", x"02",
    x"cb", x"d4", x"de", x"0c", x"10", x"7e", x"07", x"eb",
    x"d9", x"fc", x"a5", x"d9", x"cd", x"c7", x"e8", x"fd",
    x"a8", x"b2", x"00", x"f5", x"e4", x"0f", x"48", x"09",
    x"d8", x"e6", x"f1", x"d6", x"71", x"db", x"ed", x"c5",
    x"11", x"13", x"72", x"e9", x"9a", x"c0", x"12", x"26",
    x"40", x"61", x"16", x"20", x"5c", x"11", x"15", x"f9",
    x"00", x"ed", x"74", x"c7", x"31", x"a7", x"b1", x"9f",
    x"0f", x"e3", x"f7", x"e9", x"32", x"e9", x"d5", x"a9",
    x"19", x"02", x"28", x"20", x"ed", x"e5", x"fc", x"05",
    x"c5", x"12", x"17", x"1a", x"43", x"e7", x"d6", x"0b",
    x"18", x"df", x"f7", x"e9", x"bb", x"04", x"c0", x"01",
    x"06", x"04", x"01", x"ff", x"03", x"00", x"fc", x"07",
    x"3d", x"01", x"af", x"a3", x"f0", x"01", x"d8", x"fa",
    x"e7", x"05", x"02", x"07", x"f9", x"fe", x"fd", x"01",
    x"07", x"fe", x"e4", x"1a", x"df", x"1d", x"f2", x"e3",
    x"c3", x"dd", x"21", x"19", x"f7", x"05", x"c0", x"c9",
    x"eb", x"e6", x"ea", x"ee", x"e5", x"01", x"26", x"f2",
    x"0f", x"0e", x"ec", x"f7", x"0e", x"08", x"1c", x"0d",
    x"b1", x"0d", x"0b", x"83", x"e0", x"25", x"e2", x"db",
    x"06", x"8c", x"bb", x"2d", x"b6", x"17", x"34", x"e2",
    x"d4", x"2b", x"d5", x"0a", x"fc", x"20", x"cd", x"0d",
    x"00", x"b9", x"36", x"30", x"34", x"13", x"22", x"02",
    x"c6", x"00", x"1e", x"04", x"18", x"16", x"f0", x"12",
    x"ec", x"b0", x"92", x"a5", x"07", x"6e", x"ce", x"0f",
    x"25", x"ec", x"f8", x"a1", x"0c", x"e9", x"ec", x"ea",
    x"07", x"f3", x"f8", x"d6", x"b6", x"f0", x"f1", x"2a",
    x"00", x"dc", x"17", x"f6", x"d9", x"9d", x"c5", x"db",
    x"c3", x"19", x"16", x"c8", x"0f", x"0f", x"0e", x"05",
    x"11", x"91", x"e7", x"f3", x"56", x"26", x"2a", x"b8",
    x"fd", x"0d", x"6f", x"46", x"13", x"09", x"39", x"15",
    x"f9", x"dd", x"d3", x"7d", x"de", x"15", x"d8", x"23",
    x"ff", x"cb", x"d0", x"df", x"e1", x"d6", x"ce", x"ce",
    x"d3", x"14", x"0e", x"e8", x"ef", x"07", x"01", x"fb",
    x"e9", x"1a", x"fa", x"f4", x"c6", x"e7", x"78", x"41",
    x"08", x"fe", x"3c", x"32", x"11", x"07", x"18", x"b2",
    x"ff", x"ed", x"b4", x"46", x"12", x"ee", x"fc", x"d5",
    x"8a", x"96", x"de", x"f6", x"e8", x"31", x"08", x"fb",
    x"0f", x"ff", x"fb", x"ee", x"e4", x"d6", x"05", x"ff",
    x"f4", x"e1", x"cc", x"29", x"bc", x"41", x"1a", x"0c",
    x"e5", x"ae", x"04", x"17", x"f4", x"3b", x"fc", x"06",
    x"0f", x"ef", x"05", x"1f", x"fe", x"24", x"f8", x"3a",
    x"17", x"05", x"0c", x"12", x"71", x"fc", x"f2", x"f7",
    x"f2", x"0d", x"6f", x"47", x"e8", x"f5", x"f2", x"31",
    x"29", x"0b", x"2d", x"36", x"e2", x"12", x"fc", x"fc",
    x"1d", x"0e", x"db", x"e8", x"f7", x"bd", x"19", x"05",
    x"00", x"df", x"ce", x"ba", x"dd", x"34", x"da", x"16",
    x"0b", x"da", x"e9", x"cc", x"02", x"19", x"22", x"02",
    x"fa", x"03", x"f9", x"01", x"fa", x"00", x"04", x"fc",
    x"ea", x"d3", x"fd", x"0f", x"f5", x"37", x"00", x"e9",
    x"bb", x"02", x"05", x"fd", x"05", x"05", x"01", x"01",
    x"06", x"00", x"ee", x"c0", x"e1", x"cf", x"17", x"e3",
    x"15", x"fc", x"f7", x"29", x"19", x"e8", x"f8", x"fd",
    x"fd", x"0b", x"36", x"97", x"da", x"d9", x"f2", x"f5",
    x"fb", x"3a", x"f5", x"e8", x"27", x"de", x"ee", x"fa",
    x"fa", x"fc", x"29", x"23", x"e0", x"cc", x"b8", x"2b",
    x"d8", x"b3", x"2c", x"eb", x"e7", x"11", x"d1", x"d8",
    x"ab", x"d6", x"0d", x"23", x"15", x"22", x"00", x"41",
    x"ee", x"f7", x"b6", x"12", x"16", x"ee", x"d4", x"f2",
    x"e9", x"f6", x"1b", x"06", x"15", x"dc", x"cd", x"e3",
    x"bb", x"eb", x"c2", x"cd", x"f8", x"e9", x"39", x"00",
    x"ba", x"0e", x"29", x"22", x"d5", x"f4", x"b5", x"10",
    x"b0", x"ca", x"26", x"cb", x"e3", x"fb", x"f5", x"10",
    x"12", x"08", x"08", x"2b", x"50", x"af", x"21", x"19",
    x"05", x"2e", x"19", x"14", x"07", x"2c", x"d0", x"dd",
    x"05", x"18", x"b6", x"0b", x"53", x"de", x"03", x"24",
    x"3b", x"2d", x"c5", x"bc", x"f5", x"ea", x"d4", x"a2",
    x"16", x"81", x"86", x"26", x"47", x"24", x"25", x"fa",
    x"5f", x"03", x"3e", x"02", x"a3", x"01", x"ed", x"e5",
    x"1f", x"c9", x"ec", x"1a", x"05", x"25", x"f6", x"ff",
    x"26", x"da", x"f8", x"19", x"09", x"bc", x"ee", x"f2",
    x"e2", x"f1", x"e7", x"fd", x"d6", x"fe", x"2c", x"1d",
    x"d2", x"ea", x"19", x"27", x"23", x"1c", x"c2", x"d9",
    x"16", x"2f", x"e5", x"2b", x"18", x"f8", x"f6", x"cb",
    x"d8", x"e4", x"98", x"f8", x"15", x"a9", x"f0", x"b2",
    x"6c", x"ec", x"2b", x"f8", x"ed", x"13", x"22", x"28",
    x"1a", x"30", x"09", x"00", x"0c", x"26", x"0e", x"eb",
    x"06", x"c5", x"07", x"f8", x"0f", x"e4", x"a3", x"09",
    x"7a", x"98", x"e8", x"3c", x"e9", x"0b", x"40", x"c3",
    x"08", x"08", x"0e", x"f0", x"1d", x"1d", x"37", x"fe",
    x"c1", x"2c", x"18", x"dd", x"00", x"a1", x"ed", x"11",
    x"d1", x"93", x"0d", x"a5", x"d0", x"f7", x"ff", x"26",
    x"09", x"0b", x"ca", x"d2", x"30", x"fe", x"1e", x"21",
    x"f7", x"1d", x"0d", x"f5", x"f2", x"0d", x"1f", x"f9",
    x"fb", x"05", x"01", x"05", x"fc", x"fc", x"03", x"fb",
    x"fa", x"df", x"a4", x"f3", x"e9", x"9c", x"0c", x"2d",
    x"dc", x"03", x"02", x"05", x"04", x"04", x"fc", x"fb",
    x"03", x"f9", x"fa", x"3e", x"e7", x"07", x"08", x"c8",
    x"08", x"8a", x"fe", x"d0", x"44", x"fe", x"f2", x"0a",
    x"06", x"f9", x"a6", x"35", x"ee", x"c8", x"c0", x"25",
    x"13", x"d3", x"37", x"11", x"e0", x"fe", x"e9", x"04",
    x"15", x"b6", x"b9", x"04", x"ce", x"e8", x"d4", x"ef",
    x"a5", x"43", x"1a", x"e7", x"10", x"0e", x"0a", x"0f",
    x"03", x"35", x"1b", x"f6", x"fc", x"4b", x"19", x"f4",
    x"f7", x"06", x"d1", x"e1", x"ce", x"7b", x"ca", x"23",
    x"dd", x"e1", x"dc", x"e3", x"02", x"90", x"d0", x"06",
    x"12", x"ea", x"ee", x"0b", x"11", x"e8", x"ff", x"fb",
    x"12", x"d5", x"e7", x"20", x"0e", x"20", x"09", x"18",
    x"88", x"1f", x"13", x"a5", x"13", x"02", x"fb", x"ef",
    x"b9", x"27", x"02", x"11", x"11", x"ec", x"f5", x"f2",
    x"36", x"1c", x"bd", x"11", x"de", x"04", x"df", x"d8",
    x"b2", x"25", x"19", x"07", x"52", x"ef", x"db", x"00",
    x"e8", x"fd", x"26", x"14", x"b8", x"e5", x"f3", x"2f",
    x"e3", x"f7", x"13", x"0a", x"89", x"81", x"fb", x"d9",
    x"98", x"01", x"fd", x"bb", x"2d", x"1a", x"bf", x"e5",
    x"c4", x"0d", x"f1", x"c6", x"b4", x"1d", x"df", x"9a",
    x"f6", x"c4", x"f0", x"03", x"e7", x"e7", x"f1", x"10",
    x"f3", x"00", x"13", x"02", x"fe", x"de", x"e5", x"35",
    x"18", x"f0", x"0c", x"e7", x"c6", x"da", x"01", x"02",
    x"0b", x"d7", x"e0", x"15", x"24", x"c0", x"f8", x"da",
    x"d8", x"ed", x"ed", x"f2", x"03", x"07", x"f2", x"1c",
    x"fd", x"2e", x"14", x"e1", x"eb", x"2c", x"2c", x"f3",
    x"00", x"e0", x"00", x"12", x"0b", x"fd", x"07", x"f4",
    x"c6", x"11", x"0d", x"ef", x"18", x"24", x"0e", x"1c",
    x"31", x"2d", x"ce", x"25", x"f3", x"f8", x"d6", x"dd",
    x"19", x"21", x"95", x"33", x"e9", x"06", x"01", x"37",
    x"02", x"dd", x"f8", x"f3", x"e2", x"06", x"52", x"fe",
    x"eb", x"cf", x"c0", x"35", x"22", x"fa", x"ff", x"ff",
    x"f2", x"c7", x"aa", x"d8", x"09", x"e7", x"dd", x"f1",
    x"82", x"f0", x"3a", x"ed", x"e8", x"fb", x"18", x"fb",
    x"ff", x"f9", x"01", x"02", x"fd", x"07", x"05", x"fb",
    x"37", x"29", x"ff", x"2c", x"35", x"46", x"e5", x"1b",
    x"04", x"06", x"f9", x"fc", x"fa", x"05", x"03", x"fb",
    x"07", x"fd", x"f6", x"fd", x"2c", x"fc", x"85", x"1b",
    x"14", x"bc", x"e3", x"5c", x"fe", x"ed", x"27", x"32",
    x"19", x"0c", x"1b", x"01", x"24", x"11", x"fc", x"10",
    x"17", x"8b", x"d8", x"df", x"b9", x"04", x"fd", x"be",
    x"f4", x"d8", x"e9", x"d6", x"01", x"08", x"d4", x"f9",
    x"1e", x"bd", x"a9", x"0e", x"99", x"d0", x"be", x"ff",
    x"f6", x"ff", x"d6", x"f0", x"e0", x"11", x"f9", x"df",
    x"12", x"de", x"10", x"fb", x"e1", x"20", x"a5", x"12",
    x"f2", x"d7", x"b8", x"e6", x"e6", x"f8", x"b6", x"d3",
    x"12", x"04", x"00", x"ec", x"99", x"08", x"e2", x"72",
    x"d0", x"0c", x"ac", x"c6", x"e0", x"10", x"09", x"f3",
    x"e9", x"d2", x"1a", x"49", x"2d", x"3b", x"cf", x"04",
    x"30", x"03", x"2d", x"f5", x"2f", x"ff", x"f3", x"19",
    x"09", x"01", x"31", x"b1", x"2c", x"20", x"fc", x"e3",
    x"fa", x"24", x"0c", x"11", x"c9", x"15", x"e8", x"f2",
    x"ff", x"e7", x"d3", x"bf", x"06", x"f3", x"14", x"c7",
    x"07", x"e1", x"f2", x"48", x"34", x"f0", x"ae", x"1d",
    x"2f", x"12", x"e2", x"99", x"0d", x"1f", x"1d", x"e9",
    x"27", x"46", x"ee", x"fc", x"eb", x"24", x"fb", x"ef",
    x"de", x"09", x"06", x"d0", x"f6", x"19", x"1f", x"fc",
    x"b3", x"f5", x"fe", x"e8", x"f2", x"f4", x"d7", x"f5",
    x"dc", x"f8", x"ca", x"c1", x"dd", x"ed", x"f5", x"d0",
    x"28", x"1b", x"e9", x"11", x"22", x"a6", x"03", x"29",
    x"07", x"e0", x"1d", x"e9", x"dd", x"0b", x"d2", x"12",
    x"04", x"02", x"f3", x"d3", x"90", x"05", x"ea", x"db",
    x"f7", x"cf", x"e0", x"a6", x"fd", x"3f", x"f4", x"ec",
    x"e5", x"1f", x"d5", x"19", x"ca", x"d4", x"37", x"db",
    x"07", x"21", x"25", x"0d", x"8f", x"00", x"03", x"96",
    x"d7", x"35", x"f9", x"e4", x"1d", x"2b", x"26", x"19",
    x"f6", x"1a", x"ca", x"16", x"fd", x"ee", x"96", x"ef",
    x"e1", x"aa", x"34", x"24", x"0f", x"28", x"0e", x"11",
    x"f0", x"04", x"03", x"1c", x"f6", x"e3", x"d1", x"b3",
    x"de", x"1b", x"3c", x"49", x"03", x"13", x"1a", x"fc",
    x"06", x"fa", x"00", x"00", x"fa", x"fa", x"04", x"01",
    x"f0", x"0e", x"30", x"eb", x"ce", x"f6", x"14", x"fd",
    x"ef", x"ff", x"06", x"04", x"f9", x"fc", x"f9", x"04",
    x"fe", x"05", x"da", x"2c", x"f0", x"ca", x"e8", x"d4",
    x"dc", x"f3", x"0e", x"d5", x"eb", x"16", x"eb", x"e5",
    x"2b", x"06", x"ce", x"3f", x"37", x"fc", x"e2", x"07",
    x"d5", x"e4", x"1e", x"16", x"3a", x"df", x"e9", x"d8",
    x"b1", x"bb", x"c2", x"03", x"fd", x"19", x"f9", x"0a",
    x"10", x"0b", x"fc", x"ff", x"15", x"01", x"21", x"00",
    x"f7", x"26", x"2d", x"ba", x"e2", x"f9", x"ff", x"04",
    x"31", x"e4", x"bb", x"ea", x"38", x"a4", x"09", x"f8",
    x"de", x"43", x"f4", x"c8", x"f1", x"ef", x"ec", x"e5",
    x"ed", x"18", x"bf", x"f0", x"e2", x"ed", x"3a", x"f4",
    x"f6", x"10", x"0f", x"92", x"e2", x"9c", x"46", x"4e",
    x"fe", x"43", x"07", x"20", x"31", x"37", x"f9", x"0e",
    x"1b", x"e6", x"f1", x"47", x"1c", x"c7", x"b9", x"e9",
    x"1c", x"09", x"2d", x"fc", x"10", x"1d", x"1f", x"12",
    x"c9", x"c9", x"d5", x"f4", x"0c", x"fb", x"05", x"03",
    x"e9", x"ee", x"f2", x"1a", x"f9", x"1f", x"fe", x"f3",
    x"f3", x"1b", x"d1", x"33", x"09", x"aa", x"31", x"41",
    x"27", x"72", x"ce", x"a7", x"de", x"f1", x"35", x"26",
    x"f5", x"19", x"0f", x"d3", x"cd", x"d0", x"83", x"8c",
    x"11", x"e4", x"00", x"f9", x"f5", x"f6", x"e6", x"26",
    x"c9", x"11", x"0b", x"29", x"31", x"18", x"c5", x"d3",
    x"f4", x"25", x"1b", x"05", x"08", x"16", x"11", x"19",
    x"f7", x"01", x"66", x"bf", x"16", x"e2", x"06", x"1c",
    x"0e", x"f1", x"f9", x"f6", x"ab", x"bc", x"da", x"01",
    x"15", x"26", x"ff", x"22", x"0b", x"f2", x"0e", x"1b",
    x"04", x"fc", x"f7", x"f6", x"fd", x"00", x"00", x"fd",
    x"06", x"f7", x"f9", x"f9", x"fa", x"02", x"02", x"fd",
    x"03", x"f9", x"fa", x"07", x"03", x"fc", x"f3", x"00",
    x"05", x"f6", x"0b", x"fe", x"04", x"03", x"f0", x"f5",
    x"03", x"fc", x"fa", x"f5", x"03", x"fc", x"fe", x"f1",
    x"f9", x"01", x"fb", x"fa", x"f7", x"f5", x"03", x"fd",
    x"02", x"f8", x"fd", x"ff", x"03", x"fd", x"fc", x"fc",
    x"f9", x"f5", x"f3", x"fc", x"00", x"ff", x"02", x"01",
    x"01", x"fe", x"00", x"04", x"04", x"02", x"06", x"01",
    x"fc", x"fc", x"05", x"ff", x"f4", x"fb", x"01", x"f7",
    x"fe", x"fb", x"fc", x"fb", x"03", x"fd", x"01", x"05",
    x"05", x"00", x"fa", x"00", x"f8", x"fb", x"02", x"fa",
    x"fb", x"fc", x"fe", x"fc", x"ff", x"f5", x"00", x"01",
    x"01", x"f5", x"fd", x"06", x"ff", x"f8", x"fa", x"fb",
    x"f0", x"00", x"ff", x"fe", x"fc", x"fb", x"fc", x"03",
    x"f5", x"f6", x"03", x"fc", x"f9", x"00", x"f9", x"fa",
    x"04", x"02", x"fb", x"fc", x"fe", x"fc", x"f8", x"fb",
    x"03", x"fe", x"fe", x"fd", x"fc", x"fa", x"07", x"fa",
    x"04", x"fb", x"fd", x"f7", x"00", x"fd", x"f7", x"f9",
    x"f9", x"05", x"f8", x"02", x"fa", x"04", x"01", x"fd",
    x"fa", x"01", x"f7", x"03", x"04", x"fe", x"fb", x"ff",
    x"fd", x"f7", x"f6", x"fa", x"f6", x"06", x"00", x"f1",
    x"fd", x"ff", x"f0", x"02", x"f7", x"fe", x"0a", x"02",
    x"fb", x"fe", x"f8", x"02", x"fb", x"f1", x"f2", x"03",
    x"fe", x"f5", x"03", x"fe", x"fb", x"00", x"00", x"f7",
    x"fd", x"02", x"fd", x"ff", x"fc", x"00", x"ff", x"00",
    x"fd", x"00", x"fe", x"f9", x"fe", x"f4", x"f5", x"fd",
    x"00", x"fc", x"fe", x"03", x"fc", x"fb", x"f9", x"f6",
    x"f5", x"f8", x"fd", x"06", x"fb", x"f8", x"04", x"ff",
    x"02", x"ff", x"f9", x"f7", x"f8", x"02", x"ff", x"fd",
    x"f6", x"fa", x"01", x"02", x"fd", x"04", x"f7", x"05",
    x"fa", x"f8", x"f8", x"fb", x"fd", x"f2", x"01", x"f2",
    x"f1", x"f7", x"f2", x"f2", x"ff", x"fb", x"00", x"f6",
    x"01", x"f9", x"00", x"fb", x"02", x"f8", x"fe", x"f0",
    x"fb", x"01", x"fb", x"05", x"f6", x"f9", x"ff", x"f4",
    x"00", x"fc", x"fd", x"f6", x"00", x"fb", x"f7", x"01",
    x"00", x"0c", x"e2", x"28", x"26", x"03", x"fb", x"19",
    x"1c", x"11", x"ec", x"ee", x"15", x"26", x"29", x"f4",
    x"07", x"29", x"26", x"00", x"36", x"c7", x"d7", x"20",
    x"b3", x"15", x"d7", x"23", x"13", x"1e", x"56", x"1c",
    x"4b", x"c8", x"e8", x"0a", x"f2", x"ba", x"04", x"e9",
    x"c6", x"09", x"20", x"0d", x"05", x"0a", x"18", x"08",
    x"f6", x"0b", x"49", x"0e", x"e7", x"d4", x"ef", x"0a",
    x"19", x"14", x"ea", x"f2", x"b6", x"99", x"ca", x"03",
    x"ff", x"f9", x"fa", x"00", x"fd", x"00", x"fd", x"fa",
    x"1e", x"07", x"01", x"1b", x"00", x"d0", x"1b", x"10",
    x"0d", x"f9", x"ff", x"ff", x"fe", x"07", x"07", x"ff",
    x"fb", x"05", x"fe", x"1f", x"e4", x"fd", x"14", x"ed",
    x"d2", x"e1", x"0a", x"ce", x"f2", x"23", x"f7", x"14",
    x"ef", x"1f", x"29", x"2e", x"ca", x"fd", x"2c", x"18",
    x"1d", x"31", x"c8", x"db", x"f0", x"fb", x"2d", x"09",
    x"49", x"5f", x"17", x"fa", x"f1", x"f6", x"01", x"60",
    x"f0", x"28", x"f1", x"20", x"37", x"dd", x"cd", x"3d",
    x"e7", x"f1", x"fb", x"d8", x"24", x"0c", x"0a", x"d1",
    x"06", x"23", x"f8", x"f4", x"42", x"4a", x"a7", x"07",
    x"b6", x"f6", x"f6", x"35", x"fa", x"d3", x"3f", x"3b",
    x"d3", x"1a", x"08", x"ed", x"0a", x"29", x"0c", x"d9",
    x"c5", x"30", x"f2", x"bf", x"0e", x"e7", x"f4", x"1b",
    x"9e", x"38", x"c7", x"a6", x"0a", x"ec", x"40", x"25",
    x"f1", x"1c", x"87", x"ce", x"20", x"18", x"3b", x"35",
    x"26", x"fb", x"06", x"f2", x"07", x"e0", x"eb", x"df",
    x"07", x"29", x"df", x"4a", x"d5", x"04", x"1a", x"14",
    x"e2", x"f6", x"bf", x"f4", x"b9", x"29", x"f0", x"dd",
    x"15", x"23", x"2e", x"15", x"0d", x"13", x"75", x"e4",
    x"fe", x"22", x"f3", x"fd", x"2b", x"16", x"d2", x"32",
    x"fa", x"0d", x"0d", x"08", x"f7", x"22", x"ea", x"33",
    x"eb", x"cb", x"fb", x"12", x"f2", x"9c", x"ed", x"c1",
    x"c8", x"ec", x"c4", x"03", x"f0", x"d8", x"04", x"0d",
    x"1f", x"48", x"03", x"28", x"f4", x"26", x"fd", x"c4",
    x"fe", x"14", x"e1", x"01", x"08", x"01", x"0c", x"f4",
    x"08", x"12", x"a5", x"bd", x"da", x"d9", x"ca", x"21",
    x"f8", x"d6", x"73", x"e3", x"05", x"e1", x"d2", x"e6",
    x"a4", x"8d", x"cf", x"0c", x"04", x"df", x"2a", x"06",
    x"8c", x"ab", x"d9", x"ed", x"e5", x"c2", x"b2", x"97",
    x"8c", x"d2", x"25", x"20", x"2e", x"3a", x"16", x"31",
    x"12", x"30", x"2c", x"fa", x"f7", x"ff", x"28", x"02",
    x"ee", x"32", x"0e", x"03", x"c0", x"fd", x"0e", x"ef",
    x"1a", x"e0", x"0a", x"e5", x"04", x"f1", x"09", x"35",
    x"10", x"e4", x"2c", x"43", x"e1", x"20", x"05", x"d9",
    x"17", x"4b", x"f9", x"e9", x"fb", x"dd", x"00", x"02",
    x"01", x"06", x"ff", x"01", x"02", x"fe", x"fa", x"02",
    x"f2", x"a5", x"c6", x"d6", x"bd", x"e3", x"ca", x"2a",
    x"e7", x"02", x"01", x"ff", x"f9", x"f9", x"02", x"02",
    x"05", x"02", x"0c", x"04", x"b7", x"df", x"cd", x"a5",
    x"d6", x"e5", x"06", x"99", x"e8", x"c5", x"ec", x"02",
    x"01", x"cf", x"f0", x"e2", x"21", x"2c", x"18", x"0c",
    x"08", x"f4", x"f3", x"2e", x"2b", x"df", x"73", x"a2",
    x"df", x"a6", x"d0", x"7e", x"08", x"56", x"fa", x"19",
    x"22", x"ed", x"19", x"38", x"df", x"03", x"f4", x"db",
    x"23", x"35", x"08", x"32", x"f0", x"50", x"09", x"e5",
    x"3e", x"35", x"0a", x"17", x"01", x"2a", x"43", x"4b",
    x"31", x"eb", x"16", x"1c", x"02", x"0e", x"0b", x"36",
    x"16", x"25", x"f0", x"fa", x"df", x"10", x"1c", x"c9",
    x"d6", x"9a", x"17", x"1e", x"e1", x"07", x"1e", x"25",
    x"e6", x"ec", x"e7", x"31", x"20", x"44", x"0d", x"24",
    x"a9", x"44", x"b8", x"f1", x"01", x"f5", x"8a", x"ed",
    x"9c", x"a5", x"c9", x"93", x"7e", x"db", x"eb", x"f9",
    x"03", x"7f", x"db", x"df", x"80", x"e0", x"03", x"bd",
    x"1b", x"1d", x"22", x"21", x"36", x"0d", x"43", x"18",
    x"e8", x"12", x"f2", x"f6", x"e6", x"03", x"f1", x"0e",
    x"11", x"f2", x"c3", x"aa", x"00", x"92", x"51", x"6c",
    x"a1", x"83", x"cc", x"e0", x"b2", x"be", x"da", x"d9",
    x"fe", x"e9", x"0d", x"19", x"0b", x"10", x"03", x"08",
    x"03", x"f2", x"ea", x"05", x"bc", x"26", x"21", x"ca",
    x"e4", x"26", x"f4", x"1a", x"09", x"d4", x"2e", x"49",
    x"36", x"33", x"e9", x"b0", x"56", x"19", x"dc", x"03",
    x"d2", x"0e", x"ed", x"c9", x"f9", x"f0", x"f2", x"f7",
    x"09", x"fb", x"1d", x"07", x"f2", x"21", x"eb", x"fd",
    x"ee", x"08", x"06", x"03", x"ee", x"1f", x"0a", x"f4",
    x"e2", x"f5", x"f5", x"e7", x"47", x"2f", x"32", x"09",
    x"e5", x"30", x"53", x"2e", x"0d", x"ec", x"01", x"dc",
    x"41", x"51", x"38", x"f7", x"ed", x"0a", x"f0", x"14",
    x"08", x"07", x"00", x"0a", x"11", x"28", x"e1", x"0d",
    x"07", x"43", x"02", x"c6", x"3a", x"15", x"15", x"2b",
    x"e7", x"d6", x"e7", x"c2", x"34", x"51", x"a0", x"ce",
    x"e7", x"fb", x"e9", x"07", x"0b", x"dc", x"1b", x"04",
    x"fa", x"04", x"00", x"02", x"ff", x"fc", x"fb", x"03",
    x"23", x"ff", x"f0", x"f9", x"07", x"01", x"bb", x"00",
    x"24", x"00", x"fa", x"fe", x"fb", x"fc", x"00", x"fd",
    x"01", x"fc", x"fe", x"18", x"e6", x"29", x"f6", x"04",
    x"3a", x"2a", x"1a", x"2b", x"11", x"fb", x"f8", x"19",
    x"42", x"ed", x"20", x"13", x"f4", x"f7", x"06", x"d3",
    x"04", x"12", x"f5", x"ed", x"1c", x"01", x"05", x"d0",
    x"10", x"07", x"36", x"88", x"67", x"3d", x"ef", x"d9",
    x"fc", x"97", x"ca", x"01", x"d7", x"ca", x"2a", x"44",
    x"0c", x"f5", x"49", x"21", x"9f", x"1e", x"f3", x"36",
    x"f0", x"12", x"0d", x"f2", x"06", x"d5", x"0c", x"35",
    x"24", x"06", x"4c", x"09", x"24", x"06", x"00", x"1c",
    x"18", x"42", x"10", x"10", x"dc", x"f3", x"29", x"df",
    x"13", x"13", x"1d", x"f4", x"f7", x"06", x"f9", x"17",
    x"dc", x"3d", x"05", x"f7", x"45", x"05", x"09", x"0f",
    x"fd", x"0b", x"f7", x"25", x"0a", x"01", x"d5", x"ce",
    x"12", x"fc", x"27", x"3d", x"11", x"2d", x"56", x"2a",
    x"06", x"d2", x"f4", x"0a", x"89", x"75", x"08", x"f3",
    x"03", x"d8", x"dc", x"05", x"14", x"e9", x"1f", x"ef",
    x"18", x"0c", x"0d", x"de", x"fe", x"35", x"fd", x"0a",
    x"60", x"db", x"e0", x"f5", x"f8", x"0f", x"28", x"30",
    x"df", x"ee", x"2f", x"02", x"9e", x"ea", x"06", x"f0",
    x"bf", x"e5", x"36", x"e4", x"fe", x"cf", x"07", x"25",
    x"19", x"27", x"d4", x"dd", x"46", x"2d", x"2c", x"a2",
    x"c0", x"fc", x"8c", x"90", x"28", x"fc", x"dd", x"00",
    x"06", x"17", x"44", x"0b", x"dc", x"07", x"f2", x"eb",
    x"d1", x"f2", x"a2", x"b2", x"da", x"d8", x"d0", x"1f",
    x"fe", x"f0", x"44", x"3a", x"a7", x"21", x"08", x"29",
    x"b9", x"9f", x"2a", x"d0", x"fd", x"e7", x"45", x"17",
    x"c7", x"b6", x"2b", x"21", x"d1", x"03", x"06", x"12",
    x"07", x"05", x"2c", x"30", x"3d", x"36", x"db", x"e7",
    x"98", x"85", x"2b", x"86", x"de", x"02", x"03", x"31",
    x"f7", x"b9", x"dc", x"0d", x"09", x"df", x"f6", x"1b",
    x"ef", x"02", x"17", x"22", x"1c", x"20", x"09", x"d0",
    x"2a", x"10", x"f5", x"b7", x"00", x"1d", x"dc", x"0e",
    x"18", x"b6", x"ef", x"f3", x"ef", x"fd", x"fa", x"fe",
    x"fb", x"fb", x"00", x"fa", x"f9", x"f9", x"03", x"05",
    x"2e", x"dc", x"ec", x"11", x"05", x"00", x"21", x"e8",
    x"c7", x"fc", x"04", x"f9", x"04", x"04", x"02", x"fa",
    x"02", x"fa", x"9e", x"fa", x"02", x"d6", x"14", x"e9",
    x"e8", x"38", x"02", x"0f", x"1b", x"12", x"bf", x"f5",
    x"f4", x"23", x"09", x"e9", x"22", x"16", x"20", x"fa",
    x"ff", x"17", x"21", x"c3", x"23", x"14", x"eb", x"0a",
    x"1c", x"16", x"f8", x"3c", x"08", x"bc", x"ad", x"2d",
    x"07", x"07", x"4f", x"0c", x"86", x"e3", x"0d", x"fc",
    x"1e", x"05", x"e6", x"ef", x"fd", x"df", x"c0", x"0f",
    x"07", x"2b", x"08", x"25", x"14", x"15", x"dc", x"33",
    x"24", x"11", x"17", x"e5", x"0e", x"0c", x"2a", x"fb",
    x"dd", x"1d", x"c8", x"10", x"1f", x"e5", x"2c", x"e5",
    x"d8", x"00", x"45", x"f7", x"be", x"dd", x"05", x"d7",
    x"fd", x"20", x"60", x"3f", x"27", x"3e", x"03", x"f3",
    x"1c", x"ea", x"c5", x"fb", x"ed", x"c2", x"ea", x"32",
    x"1d", x"0a", x"f1", x"58", x"22", x"f5", x"dc", x"9e",
    x"e5", x"ce", x"0c", x"0a", x"68", x"03", x"26", x"04",
    x"36", x"09", x"15", x"1b", x"0d", x"0f", x"ce", x"f8",
    x"cb", x"28", x"2e", x"25", x"22", x"3d", x"16", x"11",
    x"35", x"e0", x"db", x"12", x"f9", x"07", x"11", x"22",
    x"41", x"01", x"e5", x"d9", x"16", x"20", x"c7", x"19",
    x"1f", x"e1", x"f3", x"13", x"0d", x"ec", x"0f", x"01",
    x"f3", x"20", x"fb", x"04", x"1a", x"e5", x"0b", x"0c",
    x"d6", x"02", x"25", x"1e", x"2c", x"b7", x"fd", x"27",
    x"d4", x"f3", x"23", x"11", x"f3", x"1b", x"e5", x"f7",
    x"ff", x"df", x"c2", x"d8", x"f7", x"8f", x"a1", x"82",
    x"2f", x"2a", x"96", x"ec", x"fb", x"d0", x"04", x"1d",
    x"0a", x"e6", x"15", x"1f", x"db", x"f4", x"24", x"e6",
    x"d7", x"f6", x"ec", x"06", x"f6", x"15", x"1b", x"03",
    x"24", x"6b", x"ef", x"2d", x"f3", x"2c", x"00", x"ff",
    x"39", x"b3", x"e1", x"f8", x"0b", x"3b", x"14", x"ff",
    x"1a", x"c3", x"e0", x"49", x"7b", x"15", x"30", x"93",
    x"f8", x"1e", x"4f", x"0c", x"f4", x"26", x"e5", x"aa",
    x"14", x"ed", x"bc", x"d9", x"ca", x"e5", x"f3", x"f8",
    x"f1", x"28", x"e3", x"11", x"8f", x"a0", x"f3", x"fc",
    x"04", x"04", x"07", x"ff", x"fe", x"07", x"06", x"fb",
    x"01", x"c4", x"f5", x"26", x"c4", x"16", x"01", x"91",
    x"14", x"06", x"00", x"01", x"fd", x"03", x"01", x"fc",
    x"fc", x"01", x"e7", x"14", x"cd", x"da", x"27", x"06",
    x"ea", x"f6", x"f9", x"09", x"00", x"e8", x"f3", x"2c",
    x"04", x"fb", x"3a", x"23", x"06", x"bd", x"27", x"c4",
    x"83", x"46", x"6f", x"64", x"3d", x"fa", x"38", x"fd",
    x"07", x"26", x"19", x"09", x"2a", x"0e", x"c8", x"e8",
    x"ea", x"c1", x"c7", x"d5", x"cd", x"e7", x"1c", x"09",
    x"04", x"fd", x"19", x"e8", x"14", x"11", x"a0", x"4a",
    x"00", x"cb", x"9a", x"09", x"e5", x"ba", x"cf", x"c8",
    x"e3", x"0a", x"e1", x"ec", x"1c", x"fc", x"c6", x"ab",
    x"b5", x"d5", x"0d", x"1d", x"2f", x"08", x"f5", x"14",
    x"19", x"f5", x"ef", x"0e", x"11", x"1e", x"d2", x"5d",
    x"2d", x"a4", x"c4", x"32", x"ff", x"fc", x"dd", x"4c",
    x"05", x"28", x"4b", x"d5", x"73", x"f3", x"1c", x"19",
    x"e1", x"32", x"31", x"64", x"25", x"f0", x"0d", x"f6",
    x"1c", x"d2", x"dc", x"23", x"a6", x"ef", x"f0", x"d7",
    x"0b", x"00", x"cf", x"f9", x"3b", x"e0", x"c9", x"31",
    x"08", x"e0", x"1a", x"dc", x"fe", x"05", x"cf", x"d1",
    x"07", x"fe", x"d1", x"d9", x"08", x"d5", x"f5", x"1f",
    x"bc", x"1a", x"ee", x"25", x"fa", x"d3", x"0d", x"04",
    x"ed", x"0d", x"f4", x"04", x"2d", x"1e", x"07", x"fb",
    x"f3", x"ec", x"00", x"d1", x"e3", x"f7", x"0f", x"00",
    x"00", x"f3", x"a6", x"46", x"c8", x"04", x"4b", x"10",
    x"03", x"42", x"37", x"ed", x"1f", x"24", x"09", x"d8",
    x"c4", x"ed", x"e5", x"e4", x"f2", x"df", x"d4", x"09",
    x"f9", x"f1", x"1d", x"f6", x"19", x"f9", x"f9", x"34",
    x"02", x"e3", x"1c", x"19", x"14", x"fa", x"00", x"04",
    x"9b", x"1f", x"f0", x"f9", x"e4", x"1e", x"05", x"e5",
    x"25", x"11", x"e1", x"17", x"37", x"02", x"e0", x"b7",
    x"1e", x"44", x"0f", x"08", x"c2", x"f7", x"11", x"0b",
    x"02", x"ec", x"02", x"bb", x"df", x"06", x"f1", x"ea",
    x"f0", x"0e", x"bd", x"ff", x"ef", x"db", x"df", x"ee",
    x"fd", x"b1", x"0f", x"f9", x"f1", x"d3", x"27", x"fc",
    x"0c", x"fa", x"fb", x"e1", x"1e", x"4e", x"36", x"03",
    x"01", x"fb", x"01", x"05", x"02", x"02", x"07", x"ff",
    x"07", x"df", x"01", x"c8", x"e2", x"09", x"dd", x"14",
    x"0e", x"fc", x"fb", x"ff", x"fc", x"02", x"04", x"04",
    x"f9", x"ff", x"f0", x"41", x"1b", x"14", x"0c", x"02",
    x"11", x"41", x"33", x"1e", x"e6", x"eb", x"28", x"e8",
    x"e2", x"39", x"1f", x"fe", x"10", x"f7", x"1f", x"02",
    x"ed", x"b9", x"22", x"13", x"e1", x"d3", x"d2", x"ed",
    x"dc", x"bf", x"c5", x"f7", x"01", x"11", x"85", x"f6",
    x"df", x"ee", x"af", x"2f", x"fb", x"10", x"0c", x"d7",
    x"d5", x"f5", x"ee", x"df", x"1e", x"a1", x"b0", x"ba",
    x"bf", x"cd", x"21", x"d5", x"d2", x"f3", x"07", x"de",
    x"e6", x"e9", x"fc", x"f1", x"be", x"dc", x"e4", x"da",
    x"11", x"06", x"27", x"0a", x"32", x"18", x"51", x"0d",
    x"f4", x"e8", x"fe", x"01", x"07", x"0d", x"e0", x"fe",
    x"1a", x"1f", x"e7", x"f8", x"de", x"db", x"2b", x"39",
    x"f1", x"0a", x"fa", x"32", x"dc", x"3d", x"16", x"35",
    x"ea", x"0e", x"c7", x"21", x"32", x"f4", x"c5", x"fb",
    x"1c", x"c0", x"bb", x"04", x"06", x"03", x"e0", x"d2",
    x"c4", x"d6", x"1a", x"fb", x"4b", x"f7", x"d8", x"c5",
    x"b8", x"bb", x"15", x"d5", x"ac", x"da", x"0b", x"f1",
    x"f2", x"24", x"e6", x"fa", x"fd", x"ef", x"f2", x"10",
    x"1e", x"e6", x"f6", x"02", x"05", x"bf", x"f9", x"f7",
    x"f4", x"ce", x"e8", x"05", x"17", x"09", x"0d", x"1a",
    x"f9", x"ef", x"09", x"ea", x"bc", x"eb", x"e2", x"fb",
    x"f7", x"04", x"da", x"fd", x"b4", x"e7", x"e6", x"25",
    x"28", x"0b", x"17", x"02", x"02", x"e9", x"1f", x"17",
    x"20", x"f6", x"e0", x"e0", x"e5", x"f3", x"fd", x"14",
    x"14", x"18", x"26", x"20", x"1a", x"0c", x"e3", x"ea",
    x"6b", x"bf", x"7a", x"ae", x"be", x"86", x"00", x"0d",
    x"ed", x"13", x"14", x"dd", x"29", x"d9", x"fc", x"f0",
    x"12", x"0c", x"e7", x"18", x"01", x"ed", x"bf", x"07",
    x"cd", x"9e", x"01", x"99", x"03", x"35", x"11", x"ea",
    x"f3", x"e7", x"d9", x"07", x"da", x"0f", x"06", x"dd",
    x"35", x"11", x"d5", x"25", x"14", x"c5", x"24", x"d2",
    x"21", x"d7", x"f3", x"0b", x"07", x"00", x"f0", x"fe",
    x"fd", x"fa", x"d6", x"f3", x"0a", x"e6", x"1d", x"fd",
    x"01", x"00", x"07", x"02", x"fc", x"06", x"fc", x"fe",
    x"43", x"02", x"fe", x"05", x"37", x"f8", x"21", x"fc",
    x"03", x"04", x"00", x"01", x"02", x"04", x"04", x"05",
    x"02", x"06", x"fe", x"e0", x"c0", x"1a", x"1a", x"20",
    x"f2", x"16", x"4d", x"f7", x"e6", x"d9", x"d4", x"0c",
    x"8e", x"d2", x"15", x"ed", x"f3", x"3d", x"33", x"0a",
    x"21", x"18", x"f3", x"24", x"de", x"35", x"35", x"fe",
    x"d5", x"2d", x"2a", x"c4", x"e8", x"d8", x"e9", x"45",
    x"fb", x"09", x"23", x"f7", x"d1", x"e7", x"e0", x"8d",
    x"8f", x"f3", x"25", x"4c", x"e3", x"b2", x"e5", x"ca",
    x"16", x"3f", x"1e", x"fe", x"f3", x"32", x"1c", x"01",
    x"15", x"04", x"2d", x"ff", x"08", x"f1", x"36", x"e2",
    x"1b", x"19", x"6f", x"0c", x"f0", x"fb", x"fc", x"a2",
    x"08", x"07", x"e6", x"49", x"f7", x"e2", x"c2", x"38",
    x"ee", x"0b", x"28", x"4c", x"cc", x"e9", x"0c", x"1f",
    x"08", x"ee", x"9a", x"fd", x"48", x"03", x"54", x"4f",
    x"39", x"0e", x"e4", x"07", x"1c", x"e0", x"b8", x"4f",
    x"32", x"42", x"1a", x"1c", x"4b", x"0e", x"03", x"1f",
    x"f9", x"28", x"3f", x"0f", x"13", x"24", x"df", x"0a",
    x"8c", x"39", x"1a", x"d5", x"34", x"4b", x"c6", x"06",
    x"3f", x"a5", x"44", x"00", x"00", x"fc", x"d5", x"21",
    x"42", x"fb", x"13", x"43", x"e6", x"de", x"fa", x"04",
    x"0d", x"0e", x"10", x"72", x"f2", x"e6", x"9a", x"df",
    x"a4", x"27", x"13", x"2a", x"b3", x"18", x"32", x"f8",
    x"20", x"0e", x"10", x"2e", x"e5", x"c4", x"da", x"65",
    x"9e", x"db", x"6f", x"d4", x"da", x"ca", x"e2", x"10",
    x"fb", x"c8", x"d9", x"b7", x"8d", x"80", x"90", x"6c",
    x"c1", x"9f", x"fd", x"ec", x"b9", x"07", x"cb", x"05",
    x"e4", x"ed", x"ed", x"f5", x"9f", x"9a", x"ff", x"10",
    x"b9", x"1b", x"6c", x"aa", x"ea", x"f4", x"df", x"c7",
    x"63", x"e8", x"d4", x"ee", x"f9", x"0a", x"d9", x"26",
    x"89", x"a5", x"77", x"12", x"c5", x"a9", x"12", x"f6",
    x"f3", x"70", x"1b", x"a8", x"2b", x"60", x"f3", x"f3",
    x"fd", x"26", x"b4", x"f6", x"09", x"db", x"d5", x"58",
    x"3a", x"e8", x"e8", x"2a", x"0c", x"d5", x"ef", x"0e",
    x"07", x"cc", x"d5", x"ea", x"10", x"d5", x"92", x"02",
    x"04", x"fb", x"fe", x"f9", x"07", x"03", x"04", x"fd",
    x"2f", x"3a", x"f6", x"dc", x"fe", x"bd", x"13", x"77",
    x"e6", x"01", x"fc", x"fa", x"04", x"fd", x"06", x"05",
    x"fb", x"ff", x"08", x"f0", x"e8", x"19", x"8c", x"1e",
    x"b8", x"61", x"23", x"13", x"40", x"1d", x"fd", x"cc",
    x"ec", x"ea", x"ad", x"41", x"a7", x"ec", x"df", x"f1",
    x"43", x"1d", x"1c", x"01", x"cd", x"f5", x"f1", x"ee",
    x"09", x"ed", x"1b", x"f4", x"cd", x"f7", x"2f", x"04",
    x"f7", x"16", x"16", x"e6", x"05", x"e1", x"bd", x"fd",
    x"b2", x"a7", x"00", x"0b", x"0d", x"4b", x"1e", x"28",
    x"b8", x"9d", x"14", x"1a", x"b0", x"45", x"3b", x"ce",
    x"d3", x"e0", x"f5", x"aa", x"ef", x"22", x"1a", x"0e",
    x"5b", x"ef", x"1d", x"b9", x"b8", x"f7", x"b7", x"0e",
    x"0f", x"07", x"eb", x"0a", x"36", x"c2", x"0d", x"fb",
    x"cd", x"04", x"07", x"78", x"21", x"fc", x"f0", x"09",
    x"b0", x"fa", x"23", x"e7", x"dd", x"14", x"1b", x"17",
    x"e7", x"c5", x"02", x"f0", x"5b", x"04", x"e7", x"0e",
    x"d7", x"d8", x"ff", x"0c", x"d6", x"da", x"dd", x"14",
    x"0b", x"0e", x"1b", x"2d", x"de", x"16", x"05", x"bf",
    x"28", x"df", x"c5", x"17", x"0a", x"05", x"09", x"e4",
    x"c9", x"13", x"f9", x"9b", x"10", x"f1", x"ff", x"02",
    x"f2", x"e7", x"10", x"31", x"d4", x"f5", x"b2", x"3b",
    x"d0", x"99", x"45", x"2f", x"f6", x"db", x"08", x"e5",
    x"c0", x"4a", x"27", x"07", x"df", x"ef", x"bf", x"e3",
    x"33", x"e5", x"09", x"12", x"e6", x"0f", x"91", x"56",
    x"eb", x"69", x"fb", x"06", x"cd", x"c0", x"d6", x"cc",
    x"f7", x"f1", x"ff", x"fc", x"24", x"fa", x"f0", x"0b",
    x"e0", x"dd", x"f5", x"d5", x"ba", x"5b", x"29", x"da",
    x"f6", x"fa", x"f7", x"03", x"04", x"02", x"f8", x"fb",
    x"03", x"02", x"fe", x"f7", x"fc", x"00", x"fa", x"f9",
    x"f5", x"f9", x"f9", x"f6", x"ee", x"00", x"f1", x"02",
    x"fe", x"03", x"ff", x"fb", x"f7", x"fb", x"fd", x"f2",
    x"f9", x"f7", x"ff", x"05", x"fd", x"fb", x"01", x"fd",
    x"fd", x"07", x"f2", x"00", x"f6", x"f9", x"fb", x"fa",
    x"fc", x"fa", x"fb", x"f3", x"fb", x"fa", x"02", x"00",
    x"ff", x"f3", x"f5", x"04", x"f6", x"00", x"fc", x"07",
    x"f9", x"04", x"04", x"02", x"ff", x"03", x"02", x"03",
    x"fb", x"02", x"06", x"00", x"f0", x"f8", x"00", x"06",
    x"00", x"03", x"03", x"02", x"fb", x"fd", x"fe", x"fe",
    x"05", x"fd", x"fd", x"f3", x"ff", x"fe", x"fc", x"09",
    x"f7", x"f7", x"08", x"f9", x"fd", x"f4", x"fb", x"02",
    x"07", x"fe", x"fa", x"f8", x"ff", x"f9", x"f4", x"fe",
    x"f3", x"f8", x"fa", x"01", x"fb", x"02", x"f8", x"03",
    x"ff", x"f7", x"05", x"f8", x"f8", x"09", x"f8", x"fb",
    x"f3", x"f2", x"f8", x"f8", x"f3", x"f1", x"f7", x"f7",
    x"f6", x"f0", x"fe", x"f2", x"fd", x"f9", x"f7", x"03",
    x"02", x"f8", x"fb", x"f4", x"ff", x"fc", x"01", x"02",
    x"fd", x"ff", x"00", x"f9", x"fa", x"fe", x"fc", x"fe",
    x"02", x"f7", x"f7", x"03", x"f8", x"01", x"f9", x"fc",
    x"00", x"f9", x"fe", x"01", x"00", x"04", x"fa", x"00",
    x"00", x"00", x"fe", x"fa", x"f1", x"03", x"fa", x"fa",
    x"0b", x"06", x"04", x"f4", x"fe", x"fd", x"ff", x"01",
    x"fa", x"fd", x"f6", x"05", x"f7", x"07", x"fe", x"02",
    x"fc", x"f0", x"fd", x"fa", x"f1", x"ec", x"02", x"f6",
    x"fe", x"07", x"04", x"04", x"fa", x"f1", x"03", x"04",
    x"fa", x"03", x"f6", x"fd", x"f8", x"f4", x"fc", x"00",
    x"07", x"fe", x"f3", x"0a", x"01", x"f1", x"05", x"02",
    x"f9", x"fd", x"f9", x"fc", x"ff", x"00", x"08", x"fd",
    x"fa", x"02", x"00", x"06", x"fa", x"01", x"00", x"ff",
    x"03", x"09", x"fd", x"00", x"02", x"f1", x"04", x"f8",
    x"f8", x"02", x"e9", x"f5", x"fd", x"fe", x"f8", x"02",
    x"f7", x"00", x"f5", x"f6", x"f8", x"fe", x"fa", x"fb",
    x"ef", x"f8", x"f6", x"f4", x"02", x"f6", x"fd", x"f4",
    x"f1", x"fc", x"02", x"fc", x"fd", x"f4", x"f5", x"fb",
    x"32", x"f9", x"15", x"23", x"f3", x"eb", x"e0", x"a2",
    x"bf", x"0a", x"04", x"24", x"1b", x"d6", x"2e", x"07",
    x"fc", x"ef", x"18", x"31", x"f0", x"d2", x"0f", x"f8",
    x"2d", x"38", x"47", x"3c", x"ef", x"47", x"1c", x"fc",
    x"f1", x"08", x"2e", x"f3", x"20", x"08", x"fd", x"25",
    x"18", x"25", x"e3", x"f1", x"3a", x"13", x"1b", x"a9",
    x"03", x"ea", x"b3", x"07", x"08", x"ff", x"c9", x"0b",
    x"03", x"fe", x"b0", x"9a", x"0b", x"dc", x"d3", x"fd",
    x"07", x"06", x"03", x"00", x"04", x"f9", x"03", x"ff",
    x"e9", x"f0", x"fe", x"e1", x"ca", x"21", x"25", x"be",
    x"99", x"fe", x"ff", x"fe", x"ff", x"ff", x"00", x"06",
    x"04", x"fd", x"17", x"20", x"db", x"1c", x"20", x"f4",
    x"4d", x"12", x"ef", x"dc", x"0f", x"1f", x"f5", x"0a",
    x"0e", x"38", x"e3", x"e7", x"11", x"0e", x"08", x"19",
    x"04", x"2a", x"09", x"fc", x"6a", x"06", x"31", x"42",
    x"20", x"ea", x"07", x"1a", x"c9", x"1a", x"49", x"4a",
    x"b5", x"19", x"35", x"dd", x"4a", x"09", x"17", x"48",
    x"07", x"dd", x"2e", x"06", x"ef", x"37", x"fb", x"55",
    x"29", x"ee", x"e3", x"06", x"0b", x"f5", x"11", x"1d",
    x"fd", x"02", x"bc", x"b5", x"18", x"16", x"2d", x"dc",
    x"3e", x"10", x"0a", x"0a", x"23", x"ea", x"bf", x"ee",
    x"ce", x"d8", x"fc", x"25", x"10", x"05", x"24", x"fb",
    x"01", x"03", x"f9", x"f9", x"23", x"d2", x"35", x"0b",
    x"bb", x"27", x"1c", x"04", x"0e", x"fd", x"12", x"57",
    x"e9", x"f4", x"42", x"04", x"af", x"2a", x"07", x"c7",
    x"29", x"fc", x"22", x"ed", x"e5", x"e8", x"00", x"09",
    x"e7", x"2d", x"e8", x"e8", x"11", x"95", x"d7", x"f5",
    x"29", x"49", x"25", x"f7", x"04", x"38", x"38", x"22",
    x"3e", x"c2", x"28", x"38", x"f0", x"cf", x"f1", x"d5",
    x"cb", x"b5", x"ee", x"0c", x"a8", x"d1", x"f6", x"11",
    x"e0", x"f2", x"50", x"04", x"3a", x"fd", x"ec", x"ee",
    x"ba", x"b4", x"0b", x"18", x"17", x"f2", x"d0", x"fe",
    x"21", x"10", x"02", x"1e", x"25", x"e1", x"03", x"0e",
    x"13", x"0c", x"41", x"de", x"d7", x"17", x"e9", x"a4",
    x"ec", x"d4", x"b7", x"fd", x"e0", x"d8", x"13", x"10",
    x"fc", x"b3", x"18", x"d2", x"c7", x"03", x"ee", x"03",
    x"34", x"0e", x"e9", x"da", x"ff", x"1f", x"e6", x"bd",
    x"23", x"0d", x"e8", x"e1", x"f7", x"c7", x"cb", x"32",
    x"1c", x"86", x"f6", x"d8", x"0b", x"13", x"3d", x"db",
    x"48", x"c9", x"34", x"43", x"1a", x"16", x"20", x"16",
    x"1a", x"42", x"0c", x"e3", x"3c", x"f4", x"da", x"38",
    x"15", x"94", x"15", x"f0", x"3f", x"e3", x"0d", x"20",
    x"0f", x"01", x"fe", x"fd", x"bc", x"64", x"09", x"fb",
    x"d5", x"de", x"e7", x"ea", x"e5", x"70", x"cc", x"ff",
    x"fc", x"04", x"05", x"fa", x"05", x"02", x"07", x"02",
    x"0f", x"34", x"20", x"c8", x"fe", x"a3", x"f9", x"1a",
    x"31", x"03", x"02", x"fd", x"f9", x"fb", x"01", x"fa",
    x"ff", x"00", x"0b", x"06", x"17", x"fa", x"e6", x"db",
    x"09", x"18", x"da", x"f8", x"d0", x"d9", x"04", x"70",
    x"a1", x"2c", x"a3", x"ba", x"12", x"37", x"00", x"0c",
    x"2a", x"09", x"4b", x"2c", x"ba", x"16", x"f6", x"e2",
    x"f5", x"ea", x"fb", x"29", x"09", x"f5", x"d4", x"14",
    x"0e", x"0b", x"1e", x"0a", x"4e", x"34", x"a8", x"29",
    x"30", x"32", x"2d", x"13", x"1b", x"f3", x"04", x"14",
    x"da", x"d9", x"ee", x"f7", x"ca", x"c7", x"0d", x"f2",
    x"4b", x"28", x"09", x"2f", x"de", x"da", x"c1", x"fb",
    x"8b", x"0f", x"18", x"f2", x"12", x"0a", x"0c", x"52",
    x"03", x"e2", x"cf", x"08", x"f9", x"0f", x"2d", x"3f",
    x"1b", x"ec", x"f0", x"79", x"15", x"f9", x"27", x"0f",
    x"f0", x"37", x"d3", x"13", x"d4", x"12", x"10", x"f7",
    x"04", x"d0", x"2f", x"33", x"dc", x"0c", x"2d", x"1a",
    x"f4", x"f6", x"03", x"d0", x"e7", x"18", x"cb", x"1b",
    x"00", x"21", x"34", x"31", x"06", x"0d", x"3e", x"27",
    x"f6", x"08", x"0f", x"27", x"3e", x"fa", x"39", x"06",
    x"fc", x"01", x"0e", x"c9", x"e5", x"f1", x"f2", x"c2",
    x"0e", x"3f", x"23", x"0a", x"c7", x"b9", x"da", x"6d",
    x"1f", x"e5", x"74", x"ef", x"1c", x"10", x"09", x"3b",
    x"09", x"25", x"1d", x"76", x"1f", x"2f", x"13", x"17",
    x"0b", x"d0", x"16", x"fa", x"b5", x"23", x"c7", x"e6",
    x"fd", x"dc", x"e6", x"e8", x"c9", x"bd", x"f0", x"f3",
    x"ee", x"d0", x"e5", x"c9", x"e6", x"dd", x"d9", x"0b",
    x"38", x"10", x"e1", x"00", x"08", x"fb", x"ce", x"e4",
    x"0f", x"2b", x"05", x"f6", x"f2", x"1f", x"95", x"f1",
    x"f4", x"02", x"06", x"10", x"0d", x"da", x"e1", x"32",
    x"1d", x"07", x"18", x"14", x"88", x"15", x"54", x"db",
    x"e5", x"0c", x"ea", x"0c", x"f6", x"ce", x"19", x"e4",
    x"e5", x"b9", x"2c", x"07", x"f8", x"22", x"07", x"d8",
    x"1f", x"df", x"f1", x"fe", x"d0", x"05", x"fa", x"13",
    x"da", x"d6", x"f8", x"1b", x"f2", x"5c", x"03", x"0a",
    x"f2", x"c6", x"f7", x"b2", x"8a", x"e0", x"66", x"00",
    x"02", x"ff", x"06", x"fe", x"07", x"00", x"01", x"fe",
    x"db", x"cd", x"0b", x"b5", x"ce", x"d9", x"b9", x"c9",
    x"af", x"01", x"fc", x"00", x"fc", x"fe", x"07", x"06",
    x"f9", x"00", x"1e", x"fe", x"dd", x"2c", x"f0", x"1a",
    x"c3", x"fc", x"fc", x"de", x"0d", x"ec", x"1b", x"0f",
    x"a9", x"d5", x"c6", x"c7", x"12", x"02", x"4b", x"d7",
    x"0f", x"17", x"d2", x"62", x"5d", x"f6", x"e4", x"f9",
    x"d7", x"13", x"ed", x"da", x"49", x"06", x"cc", x"c8",
    x"1f", x"da", x"25", x"1f", x"64", x"13", x"01", x"fa",
    x"14", x"12", x"cd", x"f2", x"2a", x"6e", x"17", x"20",
    x"ed", x"18", x"f1", x"dc", x"c1", x"f6", x"05", x"e2",
    x"1b", x"fb", x"f6", x"47", x"e7", x"0a", x"f3", x"1d",
    x"13", x"6a", x"1a", x"0d", x"05", x"0c", x"08", x"ef",
    x"23", x"0e", x"f2", x"0e", x"0e", x"10", x"e7", x"28",
    x"e9", x"b5", x"fd", x"d8", x"19", x"cb", x"e2", x"aa",
    x"eb", x"ad", x"86", x"30", x"79", x"0d", x"e4", x"f5",
    x"cd", x"e2", x"ee", x"36", x"51", x"10", x"1a", x"15",
    x"22", x"b9", x"04", x"08", x"39", x"40", x"15", x"88",
    x"13", x"fc", x"51", x"1b", x"46", x"46", x"1f", x"ea",
    x"0d", x"fb", x"16", x"1e", x"20", x"d1", x"2d", x"38",
    x"b0", x"02", x"eb", x"06", x"e7", x"d0", x"31", x"da",
    x"20", x"27", x"17", x"ee", x"f9", x"df", x"0c", x"ba",
    x"23", x"53", x"7f", x"09", x"0f", x"29", x"f2", x"12",
    x"25", x"96", x"f5", x"db", x"13", x"2b", x"31", x"ee",
    x"0f", x"f8", x"fe", x"11", x"f3", x"03", x"23", x"c7",
    x"07", x"e0", x"e0", x"e8", x"fd", x"eb", x"fa", x"e3",
    x"d4", x"dc", x"11", x"d6", x"c0", x"0e", x"d0", x"29",
    x"df", x"f3", x"ff", x"d5", x"f6", x"fb", x"ef", x"fe",
    x"fd", x"00", x"03", x"01", x"02", x"03", x"fd", x"01",
    x"00", x"f4", x"fa", x"fe", x"02", x"fa", x"fc", x"f8",
    x"f7", x"05", x"fe", x"ff", x"03", x"04", x"f8", x"02",
    x"01", x"fc", x"fb", x"00", x"fc", x"00", x"01", x"f9",
    x"02", x"ff", x"fa", x"01", x"fa", x"f9", x"05", x"02",
    x"f6", x"01", x"00", x"fa", x"fd", x"05", x"f8", x"fa",
    x"f4", x"fc", x"02", x"f9", x"fb", x"f7", x"f9", x"fa",
    x"fb", x"fa", x"ff", x"fa", x"00", x"f4", x"f9", x"06",
    x"fc", x"fd", x"ff", x"fe", x"02", x"ff", x"fe", x"04",
    x"f5", x"02", x"04", x"f8", x"fb", x"01", x"f9", x"f5",
    x"fa", x"06", x"06", x"04", x"01", x"fd", x"06", x"06",
    x"fb", x"fe", x"fa", x"f7", x"f7", x"f5", x"04", x"f5",
    x"fc", x"01", x"fa", x"01", x"f7", x"00", x"f8", x"f5",
    x"f8", x"00", x"01", x"f9", x"fe", x"f9", x"fd", x"fe",
    x"fc", x"fe", x"03", x"02", x"fc", x"06", x"fe", x"f9",
    x"ff", x"f7", x"ff", x"03", x"f7", x"fe", x"04", x"fa",
    x"f9", x"ff", x"06", x"ff", x"fe", x"f7", x"00", x"fb",
    x"fb", x"fe", x"fb", x"f8", x"04", x"09", x"00", x"02",
    x"f7", x"f6", x"fa", x"fb", x"ff", x"fb", x"04", x"fd",
    x"f9", x"ff", x"fa", x"fe", x"fd", x"00", x"fd", x"02",
    x"f9", x"f8", x"fb", x"fa", x"fa", x"01", x"fe", x"f4",
    x"fe", x"f6", x"01", x"fd", x"f6", x"05", x"03", x"fb",
    x"fa", x"03", x"fb", x"ff", x"04", x"01", x"01", x"ff",
    x"fe", x"f5", x"fb", x"fe", x"fc", x"00", x"00", x"ff",
    x"fa", x"f6", x"f3", x"fc", x"f7", x"ff", x"fb", x"fa",
    x"f7", x"f4", x"01", x"f3", x"05", x"f9", x"05", x"fa",
    x"fc", x"06", x"fe", x"fc", x"f6", x"01", x"f9", x"f6",
    x"01", x"fc", x"fc", x"ff", x"fd", x"ff", x"f8", x"fd",
    x"02", x"ff", x"02", x"fa", x"fc", x"fd", x"f7", x"f8",
    x"f7", x"f8", x"fc", x"01", x"fd", x"fb", x"ff", x"f8",
    x"f8", x"fd", x"fb", x"04", x"f8", x"02", x"03", x"f8",
    x"01", x"f8", x"f8", x"fc", x"f7", x"fa", x"fc", x"fb",
    x"fa", x"f8", x"fa", x"00", x"f7", x"fb", x"f7", x"ff",
    x"fb", x"01", x"fa", x"fd", x"f5", x"01", x"00", x"ff",
    x"f5", x"f5", x"f5", x"f1", x"fb", x"fc", x"f5", x"f7",
    x"fb", x"f4", x"f6", x"fd", x"f9", x"f8", x"f4", x"f3",
    x"0d", x"03", x"3a", x"f4", x"04", x"e3", x"e3", x"03",
    x"fe", x"07", x"fc", x"21", x"37", x"0c", x"32", x"29",
    x"40", x"0e", x"fc", x"d2", x"f4", x"04", x"1b", x"e9",
    x"12", x"f8", x"9d", x"f9", x"1b", x"10", x"25", x"2b",
    x"3c", x"ca", x"1c", x"45", x"9a", x"dd", x"c4", x"09",
    x"26", x"22", x"2c", x"f7", x"d8", x"f3", x"c6", x"8e",
    x"fc", x"fa", x"f0", x"c9", x"4f", x"2c", x"09", x"07",
    x"f0", x"0c", x"e4", x"b4", x"09", x"ea", x"e2", x"02",
    x"fa", x"05", x"06", x"fc", x"fc", x"06", x"07", x"06",
    x"ef", x"07", x"0b", x"ea", x"17", x"ee", x"94", x"fc",
    x"3b", x"fb", x"fa", x"06", x"fa", x"fd", x"01", x"04",
    x"00", x"02", x"ae", x"bc", x"ca", x"06", x"3e", x"0d",
    x"fd", x"e9", x"0e", x"ca", x"e7", x"cc", x"3a", x"3d",
    x"ec", x"fb", x"b9", x"bd", x"08", x"37", x"01", x"e5",
    x"ef", x"2b", x"15", x"03", x"05", x"08", x"03", x"fe",
    x"cf", x"0a", x"2b", x"e4", x"1a", x"e5", x"cb", x"d5",
    x"b9", x"21", x"af", x"f0", x"02", x"d9", x"00", x"ff",
    x"f5", x"23", x"2c", x"24", x"f8", x"cf", x"1d", x"15",
    x"18", x"cb", x"c3", x"f4", x"e5", x"d7", x"33", x"1e",
    x"83", x"e5", x"a3", x"c5", x"14", x"fc", x"3e", x"15",
    x"d6", x"b9", x"1d", x"26", x"1b", x"16", x"06", x"dc",
    x"1e", x"03", x"ed", x"0b", x"00", x"b2", x"de", x"34",
    x"2f", x"2a", x"01", x"e4", x"1a", x"fa", x"fa", x"0e",
    x"bc", x"de", x"2c", x"23", x"27", x"20", x"20", x"11",
    x"dc", x"03", x"3e", x"52", x"33", x"00", x"01", x"cb",
    x"d2", x"b4", x"b3", x"21", x"e7", x"01", x"1f", x"e7",
    x"f5", x"f5", x"ba", x"fe", x"ed", x"d6", x"2d", x"3f",
    x"d2", x"26", x"07", x"12", x"0c", x"2d", x"ed", x"11",
    x"eb", x"13", x"1b", x"06", x"27", x"19", x"03", x"1b",
    x"00", x"1f", x"f0", x"01", x"ec", x"de", x"06", x"6a",
    x"05", x"b8", x"6b", x"e0", x"e9", x"ca", x"07", x"d3",
    x"24", x"c5", x"46", x"08", x"fd", x"a2", x"b7", x"d4",
    x"ec", x"25", x"b4", x"38", x"32", x"0f", x"d6", x"f4",
    x"31", x"33", x"2e", x"02", x"e2", x"fe", x"06", x"0d",
    x"ef", x"c5", x"ed", x"f9", x"da", x"9e", x"d5", x"fc",
    x"8d", x"32", x"23", x"8d", x"f4", x"e4", x"0d", x"0d",
    x"6c", x"ed", x"13", x"bc", x"af", x"c6", x"04", x"04",
    x"15", x"bd", x"ec", x"5a", x"de", x"18", x"19", x"2e",
    x"ea", x"c2", x"0f", x"38", x"3a", x"07", x"ca", x"39",
    x"dd", x"2b", x"e7", x"ef", x"e3", x"2d", x"33", x"37",
    x"2a", x"e0", x"ff", x"fc", x"17", x"e1", x"04", x"10",
    x"1e", x"0f", x"12", x"18", x"0f", x"30", x"1b", x"b8",
    x"05", x"b7", x"fd", x"ac", x"e4", x"1f", x"0f", x"37",
    x"25", x"cf", x"dd", x"c9", x"1f", x"1d", x"76", x"04",
    x"02", x"01", x"fb", x"fc", x"fe", x"f9", x"02", x"05",
    x"d2", x"f5", x"f8", x"40", x"43", x"cc", x"0b", x"e0",
    x"9a", x"02", x"03", x"07", x"fb", x"f9", x"fa", x"02",
    x"fa", x"f9", x"e5", x"c4", x"04", x"24", x"1b", x"f6",
    x"17", x"db", x"b2", x"a3", x"e4", x"27", x"dd", x"f1",
    x"e1", x"d8", x"2a", x"42", x"f1", x"d8", x"d1", x"0b",
    x"29", x"22", x"f2", x"22", x"10", x"e2", x"c0", x"1c",
    x"d2", x"fc", x"f7", x"cb", x"f3", x"06", x"48", x"0e",
    x"c4", x"16", x"f3", x"0d", x"d2", x"19", x"20", x"1a",
    x"ea", x"d0", x"16", x"bf", x"e7", x"be", x"53", x"26",
    x"2b", x"48", x"0d", x"11", x"0a", x"1c", x"f1", x"ee",
    x"bf", x"15", x"01", x"a8", x"0c", x"eb", x"ec", x"e2",
    x"d7", x"db", x"17", x"36", x"48", x"d1", x"18", x"e9",
    x"14", x"58", x"e8", x"f6", x"e1", x"09", x"06", x"07",
    x"10", x"4f", x"3a", x"63", x"33", x"38", x"04", x"f5",
    x"06", x"21", x"ef", x"02", x"df", x"72", x"1c", x"3d",
    x"9d", x"2d", x"24", x"3e", x"27", x"cb", x"0e", x"90",
    x"e6", x"da", x"c4", x"fa", x"10", x"00", x"07", x"cd",
    x"09", x"1a", x"f9", x"fb", x"16", x"d7", x"1b", x"3b",
    x"1f", x"1e", x"11", x"25", x"07", x"dd", x"c8", x"c7",
    x"fe", x"ed", x"1d", x"58", x"08", x"0d", x"09", x"00",
    x"10", x"c4", x"fd", x"91", x"ae", x"0c", x"e4", x"d2",
    x"e7", x"c1", x"f9", x"1d", x"11", x"f0", x"07", x"e3",
    x"16", x"1a", x"1a", x"f4", x"e9", x"85", x"ab", x"09",
    x"b6", x"e9", x"fb", x"fd", x"20", x"e2", x"ff", x"48",
    x"fb", x"04", x"1a", x"24", x"59", x"10", x"ec", x"c2",
    x"e2", x"f0", x"a2", x"f7", x"f6", x"c1", x"ec", x"26",
    x"23", x"f5", x"b8", x"ff", x"fe", x"f6", x"2d", x"eb",
    x"c5", x"c5", x"f7", x"08", x"02", x"b8", x"fb", x"c8",
    x"b9", x"18", x"23", x"29", x"f0", x"e7", x"94", x"22",
    x"e4", x"a0", x"12", x"dc", x"01", x"1f", x"ee", x"5a",
    x"3a", x"4d", x"7b", x"18", x"0c", x"2f", x"4c", x"09",
    x"e8", x"fc", x"3b", x"21", x"f9", x"ea", x"6f", x"19",
    x"f9", x"0e", x"01", x"00", x"18", x"fb", x"0b", x"12",
    x"15", x"0c", x"64", x"ea", x"38", x"f1", x"fb", x"f7",
    x"a1", x"b1", x"0b", x"05", x"e4", x"f8", x"f6", x"fc",
    x"02", x"ff", x"06", x"fd", x"03", x"ff", x"02", x"fe",
    x"19", x"18", x"da", x"eb", x"24", x"37", x"ee", x"e3",
    x"e1", x"00", x"ff", x"06", x"03", x"05", x"02", x"fa",
    x"02", x"07", x"fe", x"f9", x"57", x"16", x"f9", x"f1",
    x"1f", x"1b", x"b7", x"f5", x"f7", x"b2", x"0c", x"f8",
    x"1a", x"e7", x"cf", x"95", x"16", x"0e", x"ae", x"1a",
    x"2e", x"21", x"06", x"23", x"16", x"17", x"e5", x"94",
    x"fc", x"10", x"fd", x"f2", x"12", x"07", x"d4", x"f4",
    x"33", x"12", x"f4", x"06", x"05", x"1d", x"39", x"15",
    x"01", x"3a", x"1a", x"e8", x"cd", x"d2", x"1e", x"06",
    x"02", x"c1", x"03", x"1f", x"00", x"27", x"3d", x"25",
    x"1d", x"12", x"d4", x"0f", x"28", x"fd", x"6e", x"09",
    x"41", x"53", x"14", x"1d", x"f7", x"17", x"09", x"a9",
    x"0e", x"39", x"b3", x"f5", x"fa", x"21", x"1f", x"f1",
    x"1c", x"01", x"1a", x"ec", x"25", x"45", x"fb", x"fa",
    x"11", x"ae", x"16", x"db", x"71", x"24", x"df", x"d0",
    x"eb", x"17", x"57", x"fd", x"05", x"14", x"16", x"fb",
    x"dd", x"d6", x"f7", x"3a", x"f1", x"fb", x"36", x"1c",
    x"13", x"2e", x"0d", x"e4", x"2f", x"f9", x"e4", x"0d",
    x"0d", x"e9", x"4a", x"3c", x"25", x"07", x"1d", x"3e",
    x"27", x"05", x"ea", x"99", x"f3", x"3a", x"02", x"09",
    x"cc", x"dc", x"01", x"b2", x"c2", x"01", x"dd", x"d4",
    x"e4", x"12", x"11", x"d4", x"b3", x"c7", x"19", x"42",
    x"b6", x"15", x"27", x"e0", x"4a", x"3c", x"07", x"d5",
    x"dc", x"21", x"b2", x"1d", x"4b", x"12", x"98", x"3e",
    x"00", x"d3", x"d4", x"06", x"04", x"06", x"f5", x"f1",
    x"f3", x"b8", x"b3", x"d4", x"d2", x"f0", x"d4", x"eb",
    x"d7", x"15", x"1a", x"e2", x"81", x"29", x"30", x"de",
    x"e8", x"07", x"3b", x"d5", x"fb", x"cf", x"e3", x"0c",
    x"1b", x"e9", x"eb", x"10", x"51", x"24", x"fc", x"a7",
    x"a2", x"d3", x"e8", x"d3", x"ed", x"fd", x"17", x"03",
    x"3c", x"37", x"d0", x"17", x"24", x"fb", x"05", x"1d",
    x"29", x"eb", x"02", x"e7", x"19", x"ff", x"35", x"32",
    x"b9", x"f3", x"c7", x"e6", x"06", x"f8", x"26", x"db",
    x"f6", x"01", x"19", x"10", x"fb", x"10", x"d7", x"03",
    x"2f", x"f0", x"bd", x"cc", x"34", x"12", x"fd", x"fd",
    x"04", x"fc", x"07", x"03", x"fe", x"00", x"00", x"02",
    x"be", x"c3", x"f6", x"d4", x"0b", x"f5", x"f5", x"0b",
    x"fd", x"03", x"04", x"ff", x"06", x"fe", x"f9", x"04",
    x"00", x"04", x"ea", x"30", x"18", x"ea", x"0e", x"09",
    x"c7", x"07", x"2c", x"81", x"0d", x"35", x"24", x"07",
    x"0a", x"f5", x"ab", x"68", x"58", x"07", x"ec", x"0f",
    x"f8", x"2b", x"fc", x"05", x"17", x"83", x"ce", x"39",
    x"d5", x"0e", x"2a", x"d2", x"cd", x"b4", x"f3", x"3d",
    x"29", x"c6", x"19", x"07", x"00", x"0e", x"cb", x"3e",
    x"29", x"03", x"02", x"08", x"11", x"10", x"1d", x"5b",
    x"29", x"0d", x"ee", x"af", x"02", x"17", x"23", x"12",
    x"be", x"57", x"1c", x"28", x"08", x"08", x"1f", x"20",
    x"19", x"eb", x"ea", x"fa", x"f8", x"f2", x"f8", x"f7",
    x"af", x"08", x"fd", x"13", x"f3", x"1a", x"12", x"b9",
    x"1a", x"22", x"d0", x"14", x"fe", x"db", x"8b", x"26",
    x"3b", x"fb", x"2f", x"36", x"dd", x"0a", x"be", x"05",
    x"c3", x"c7", x"07", x"22", x"1e", x"31", x"c4", x"09",
    x"13", x"cd", x"f4", x"e5", x"6a", x"b6", x"04", x"2a",
    x"54", x"d8", x"12", x"0b", x"f1", x"d6", x"ed", x"fd",
    x"46", x"2c", x"4b", x"ec", x"ff", x"3e", x"06", x"04",
    x"2b", x"84", x"d7", x"34", x"5f", x"60", x"8a", x"cc",
    x"12", x"31", x"17", x"00", x"10", x"f5", x"db", x"17",
    x"d0", x"b0", x"bd", x"db", x"00", x"2b", x"13", x"c6",
    x"d8", x"01", x"3b", x"02", x"09", x"e3", x"e1", x"e1",
    x"dc", x"2b", x"d0", x"0a", x"2f", x"f5", x"2f", x"42",
    x"23", x"df", x"13", x"10", x"c6", x"05", x"00", x"cf",
    x"df", x"e4", x"cf", x"0f", x"e0", x"ec", x"e2", x"27",
    x"18", x"05", x"fc", x"f6", x"0d", x"e3", x"f6", x"fb",
    x"df", x"c1", x"0c", x"7c", x"0d", x"00", x"5a", x"d4",
    x"ed", x"f2", x"0f", x"2d", x"f3", x"06", x"e9", x"eb",
    x"18", x"fe", x"11", x"1d", x"01", x"24", x"1b", x"19",
    x"33", x"eb", x"2a", x"82", x"f5", x"31", x"7b", x"ed",
    x"18", x"c6", x"1f", x"1a", x"d0", x"e4", x"06", x"e7",
    x"e2", x"f1", x"02", x"33", x"dc", x"f2", x"2b", x"29",
    x"f5", x"ea", x"f3", x"f0", x"e4", x"0f", x"e5", x"d6",
    x"fb", x"c8", x"e9", x"f7", x"04", x"31", x"e8", x"01",
    x"fb", x"05", x"fc", x"fe", x"05", x"06", x"ff", x"07",
    x"e0", x"04", x"f1", x"04", x"38", x"e7", x"e2", x"d2",
    x"e8", x"05", x"03", x"04", x"ff", x"01", x"04", x"00",
    x"f9", x"fb", x"d3", x"12", x"26", x"db", x"46", x"38",
    x"04", x"00", x"06", x"ee", x"fc", x"33", x"be", x"08",
    x"2e", x"22", x"18", x"e6", x"fc", x"0d", x"e7", x"ef",
    x"36", x"e1", x"1b", x"33", x"19", x"d7", x"ff", x"33",
    x"d9", x"22", x"0c", x"3e", x"3c", x"f8", x"17", x"31",
    x"0a", x"b1", x"16", x"02", x"d1", x"ff", x"ff", x"c5",
    x"e2", x"5a", x"89", x"0b", x"1c", x"9a", x"e4", x"0b",
    x"f3", x"27", x"1c", x"07", x"e2", x"df", x"23", x"02",
    x"0d", x"f7", x"39", x"00", x"28", x"f9", x"f0", x"1f",
    x"f0", x"f1", x"73", x"26", x"34", x"c1", x"eb", x"2b",
    x"e6", x"f5", x"31", x"d1", x"00", x"c7", x"c2", x"f5",
    x"20", x"2a", x"20", x"e3", x"22", x"ec", x"05", x"ae",
    x"21", x"12", x"18", x"4b", x"ba", x"c7", x"f2", x"3b",
    x"13", x"0f", x"19", x"f3", x"45", x"0e", x"36", x"b7",
    x"fe", x"a3", x"2a", x"0d", x"ae", x"f4", x"fa", x"a8",
    x"f6", x"33", x"fd", x"0f", x"1a", x"f8", x"fc", x"0f",
    x"ad", x"fb", x"08", x"06", x"29", x"e0", x"05", x"2f",
    x"13", x"05", x"fd", x"13", x"b3", x"fd", x"ea", x"e4",
    x"2a", x"2b", x"e7", x"1b", x"2e", x"db", x"30", x"dc",
    x"ef", x"ef", x"ad", x"cd", x"07", x"f5", x"98", x"f3",
    x"c0", x"f0", x"02", x"c2", x"e6", x"3f", x"e6", x"36",
    x"28", x"f0", x"e4", x"f4", x"1e", x"e6", x"e6", x"58",
    x"01", x"fc", x"07", x"ee", x"2a", x"13", x"ef", x"f1",
    x"d1", x"da", x"e4", x"c5", x"f4", x"d8", x"de", x"58",
    x"0f", x"21", x"8e", x"06", x"21", x"78", x"cb", x"c3",
    x"0a", x"cd", x"1e", x"25", x"fd", x"1b", x"fb", x"de",
    x"d6", x"da", x"1a", x"27", x"04", x"f1", x"c6", x"64",
    x"d6", x"09", x"03", x"16", x"01", x"f7", x"f8", x"cb",
    x"7f", x"83", x"cd", x"1a", x"20", x"59", x"27", x"1b",
    x"2b", x"b9", x"ce", x"de", x"c7", x"0c", x"0d", x"25",
    x"2b", x"1a", x"fd", x"81", x"a2", x"03", x"0d", x"3b",
    x"f1", x"1d", x"0e", x"b0", x"52", x"2f", x"0e", x"f9",
    x"12", x"04", x"be", x"bf", x"7b", x"57", x"a7", x"02",
    x"02", x"00", x"02", x"04", x"fd", x"03", x"00", x"f9",
    x"d5", x"d3", x"12", x"e7", x"b3", x"17", x"b8", x"6d",
    x"10", x"ff", x"fa", x"fe", x"07", x"fb", x"fc", x"01",
    x"03", x"07", x"f5", x"e2", x"17", x"f7", x"e0", x"fc",
    x"e7", x"c3", x"da", x"38", x"dc", x"ab", x"e7", x"dd",
    x"fd", x"12", x"e9", x"bf", x"e0", x"00", x"fc", x"23",
    x"2c", x"ee", x"e4", x"c9", x"dc", x"ee", x"19", x"e4",
    x"28", x"0b", x"e2", x"df", x"dd", x"82", x"f7", x"08",
    x"36", x"f8", x"1e", x"35", x"b2", x"61", x"8e", x"07",
    x"21", x"41", x"3b", x"21", x"fe", x"0d", x"f7", x"e2",
    x"d0", x"ed", x"09", x"ec", x"f0", x"46", x"5c", x"b9",
    x"c8", x"ee", x"27", x"07", x"08", x"d7", x"da", x"af",
    x"17", x"a9", x"f5", x"2e", x"1e", x"2e", x"04", x"c5",
    x"97", x"91", x"09", x"00", x"ec", x"05", x"2b", x"1b",
    x"f9", x"3d", x"f6", x"b1", x"e0", x"fd", x"27", x"f5",
    x"e7", x"36", x"df", x"54", x"4b", x"fc", x"fa", x"03",
    x"fc", x"e3", x"a5", x"cf", x"9b", x"86", x"ec", x"e8",
    x"d6", x"df", x"fd", x"dd", x"e9", x"e9", x"ba", x"f1",
    x"16", x"44", x"1c", x"18", x"fc", x"ef", x"c1", x"59",
    x"0f", x"0e", x"20", x"0d", x"1c", x"fd", x"b5", x"bb",
    x"13", x"12", x"f0", x"27", x"fa", x"e4", x"c8", x"7a",
    x"75", x"73", x"f3", x"f5", x"e6", x"07", x"24", x"b1",
    x"0b", x"d1", x"d4", x"ef", x"ff", x"ee", x"f8", x"06",
    x"2d", x"ef", x"a1", x"d2", x"05", x"0a", x"33", x"f7",
    x"18", x"07", x"cc", x"d5", x"c6", x"11", x"f9", x"2c",
    x"19", x"ec", x"df", x"fb", x"c4", x"04", x"df", x"05",
    x"f6", x"06", x"09", x"ed", x"fe", x"05", x"fe", x"32",
    x"0b", x"2a", x"38", x"fd", x"00", x"eb", x"ed", x"0a",
    x"21", x"96", x"e3", x"fe", x"07", x"d2", x"ce", x"0b",
    x"f3", x"0e", x"e3", x"0b", x"ab", x"1d", x"16", x"3f",
    x"fa", x"1f", x"e6", x"f8", x"02", x"ce", x"d4", x"f6",
    x"c6", x"fb", x"36", x"12", x"19", x"f7", x"29", x"52",
    x"3a", x"1d", x"fe", x"35", x"e6", x"1b", x"fc", x"22",
    x"3d", x"2e", x"c3", x"a0", x"f9", x"d7", x"f1", x"c4",
    x"dc", x"fd", x"1c", x"98", x"e7", x"21", x"fe", x"29",
    x"4b", x"e1", x"e6", x"d5", x"a1", x"be", x"9d", x"03",
    x"04", x"03", x"05", x"fc", x"fe", x"fe", x"02", x"f9",
    x"27", x"e2", x"15", x"a5", x"e4", x"ba", x"1d", x"fd",
    x"b9", x"04", x"05", x"fe", x"fa", x"01", x"fe", x"fd",
    x"03", x"05", x"11", x"0f", x"25", x"56", x"eb", x"1d",
    x"f4", x"c6", x"79", x"b3", x"53", x"a3", x"d3", x"37",
    x"06", x"14", x"c0", x"b0", x"0d", x"f9", x"12", x"0a",
    x"15", x"05", x"15", x"1c", x"36", x"0a", x"b0", x"dc",
    x"e3", x"d8", x"f6", x"fb", x"ff", x"13", x"01", x"fb",
    x"07", x"41", x"f5", x"60", x"19", x"bd", x"cb", x"e8",
    x"f4", x"c6", x"3f", x"1b", x"0a", x"02", x"23", x"2d",
    x"ca", x"00", x"c4", x"c2", x"d3", x"ed", x"c3", x"f2",
    x"34", x"2b", x"fe", x"ef", x"1f", x"1e", x"25", x"fc",
    x"e1", x"0d", x"31", x"0e", x"12", x"13", x"12", x"cc",
    x"19", x"f7", x"d9", x"e8", x"12", x"29", x"1a", x"03",
    x"20", x"c3", x"df", x"ab", x"19", x"20", x"29", x"a1",
    x"82", x"d5", x"f7", x"e9", x"c4", x"0b", x"24", x"0d",
    x"04", x"13", x"b6", x"da", x"c5", x"d1", x"24", x"f3",
    x"04", x"ee", x"03", x"f7", x"31", x"f0", x"11", x"21",
    x"2b", x"e4", x"46", x"5c", x"17", x"01", x"57", x"ca",
    x"0a", x"ac", x"e9", x"f9", x"28", x"19", x"bd", x"e9",
    x"f2", x"c1", x"01", x"11", x"ea", x"2e", x"f6", x"0d",
    x"d6", x"c5", x"05", x"fa", x"fe", x"e3", x"2d", x"20",
    x"f3", x"fb", x"f6", x"1d", x"c7", x"74", x"fb", x"b3",
    x"fb", x"9f", x"d4", x"99", x"fa", x"f0", x"e8", x"e9",
    x"13", x"2a", x"e6", x"09", x"16", x"e9", x"f0", x"7a",
    x"08", x"0d", x"f7", x"02", x"eb", x"ef", x"03", x"f7",
    x"04", x"dc", x"d4", x"e6", x"e3", x"01", x"e7", x"ef",
    x"eb", x"dc", x"52", x"ed", x"11", x"b5", x"f9", x"28",
    x"f7", x"fb", x"04", x"fa", x"fb", x"f8", x"fa", x"f8",
    x"f5", x"fe", x"fa", x"ff", x"00", x"f3", x"f8", x"f8",
    x"f3", x"ff", x"01", x"f6", x"f8", x"ff", x"06", x"f7",
    x"fc", x"04", x"02", x"fc", x"02", x"f9", x"f9", x"f8",
    x"fc", x"00", x"ff", x"fb", x"ff", x"06", x"05", x"f9",
    x"f4", x"f5", x"fa", x"f8", x"02", x"f6", x"04", x"02",
    x"f8", x"01", x"ff", x"fa", x"09", x"02", x"f5", x"f0",
    x"f6", x"f8", x"f9", x"01", x"03", x"00", x"01", x"fa",
    x"fd", x"f9", x"02", x"fe", x"00", x"f9", x"03", x"05",
    x"fd", x"fb", x"04", x"00", x"fe", x"01", x"f8", x"01",
    x"04", x"fe", x"fd", x"02", x"00", x"fd", x"fd", x"02",
    x"fa", x"fc", x"01", x"ff", x"08", x"f7", x"f8", x"fa",
    x"fe", x"f7", x"fb", x"fb", x"08", x"fd", x"01", x"fa",
    x"fd", x"fe", x"ff", x"05", x"04", x"f9", x"fe", x"f8",
    x"03", x"fc", x"03", x"fd", x"f8", x"f9", x"f3", x"f5",
    x"ff", x"fe", x"fb", x"fa", x"fc", x"00", x"f6", x"06",
    x"fc", x"02", x"03", x"fc", x"f6", x"01", x"01", x"ff",
    x"04", x"02", x"fa", x"fe", x"fc", x"fc", x"fe", x"f5",
    x"fc", x"fe", x"fa", x"00", x"fa", x"f6", x"fe", x"f5",
    x"02", x"f7", x"05", x"fb", x"fd", x"f5", x"f6", x"00",
    x"f6", x"ff", x"02", x"fb", x"fe", x"fa", x"fa", x"f5",
    x"fa", x"03", x"fc", x"f6", x"04", x"02", x"fa", x"00",
    x"04", x"f6", x"00", x"fb", x"04", x"f4", x"02", x"06",
    x"07", x"f9", x"ff", x"f9", x"f7", x"00", x"01", x"f8",
    x"f9", x"fa", x"fc", x"fc", x"01", x"f5", x"fc", x"00",
    x"ff", x"f7", x"03", x"f7", x"fe", x"fc", x"f8", x"fe",
    x"fa", x"ff", x"fa", x"00", x"f9", x"fa", x"03", x"fa",
    x"ff", x"fc", x"00", x"ff", x"f7", x"f7", x"f5", x"01",
    x"fa", x"fe", x"fb", x"07", x"fa", x"f5", x"01", x"02",
    x"fe", x"fd", x"fd", x"f6", x"f9", x"02", x"fa", x"f5",
    x"04", x"f6", x"f7", x"f7", x"fa", x"fc", x"02", x"fa",
    x"fe", x"fa", x"ff", x"ff", x"f6", x"f5", x"f9", x"f7",
    x"fa", x"f3", x"f5", x"f5", x"f9", x"01", x"fe", x"07",
    x"02", x"fc", x"02", x"03", x"f5", x"fc", x"f6", x"00",
    x"fb", x"01", x"fe", x"f6", x"fd", x"f7", x"f4", x"fb",
    x"f7", x"f5", x"f8", x"f8", x"f3", x"05", x"fd", x"f9",
    x"01", x"fc", x"fb", x"f6", x"04", x"ff", x"01", x"f5",
    x"f8", x"f5", x"fe", x"fc", x"f5", x"f5", x"fd", x"fc",
    x"fc", x"f9", x"03", x"00", x"03", x"fe", x"03", x"f5",
    x"fc", x"f9", x"00", x"03", x"00", x"fd", x"fd", x"fc",
    x"03", x"fc", x"f7", x"ff", x"fe", x"fb", x"fc", x"01",
    x"02", x"f6", x"03", x"f6", x"fb", x"04", x"06", x"04",
    x"fe", x"fb", x"01", x"05", x"02", x"fb", x"f9", x"03",
    x"fe", x"f9", x"f7", x"f8", x"ff", x"f8", x"00", x"06",
    x"fb", x"01", x"fc", x"04", x"f9", x"fb", x"fb", x"03",
    x"f9", x"fb", x"02", x"fc", x"03", x"f7", x"03", x"01",
    x"f5", x"f9", x"fb", x"fe", x"05", x"05", x"07", x"f9",
    x"fa", x"07", x"fe", x"fc", x"00", x"fb", x"02", x"01",
    x"f7", x"f8", x"fd", x"fd", x"00", x"05", x"fa", x"fa",
    x"04", x"05", x"03", x"fa", x"f8", x"04", x"06", x"00",
    x"f8", x"f5", x"04", x"f9", x"00", x"01", x"f6", x"00",
    x"f7", x"fb", x"f4", x"05", x"f5", x"00", x"fd", x"f7",
    x"f6", x"fa", x"fd", x"00", x"f7", x"ff", x"04", x"fc",
    x"03", x"fb", x"ff", x"07", x"f8", x"01", x"fc", x"f9",
    x"f9", x"03", x"04", x"fb", x"03", x"03", x"fd", x"01",
    x"fd", x"01", x"fb", x"05", x"fa", x"f6", x"fe", x"fe",
    x"01", x"f9", x"02", x"fb", x"fe", x"ff", x"05", x"fc",
    x"f7", x"f7", x"f6", x"ff", x"04", x"fc", x"fd", x"00",
    x"ff", x"f6", x"ff", x"04", x"fe", x"04", x"fa", x"f7",
    x"f6", x"f7", x"ff", x"fc", x"fd", x"00", x"01", x"fb",
    x"f9", x"f5", x"f8", x"fd", x"00", x"fc", x"02", x"fb",
    x"fe", x"f8", x"fb", x"fb", x"03", x"01", x"f8", x"fc",
    x"02", x"fa", x"fa", x"f6", x"fd", x"ff", x"05", x"00",
    x"f5", x"f9", x"01", x"fb", x"f7", x"fa", x"fa", x"fc",
    x"fd", x"f5", x"01", x"f7", x"00", x"fe", x"fb", x"02",
    x"fd", x"ff", x"00", x"00", x"fb", x"f5", x"f6", x"f7",
    x"00", x"fe", x"fc", x"f7", x"fb", x"ff", x"f9", x"fc",
    x"fa", x"01", x"f8", x"fc", x"fc", x"fd", x"f6", x"fc",
    x"fd", x"f7", x"02", x"fa", x"fb", x"04", x"f6", x"03",
    x"f8", x"f7", x"02", x"fd", x"00", x"f9", x"fa", x"00",
    x"f7", x"fb", x"ff", x"fb", x"02", x"fc", x"fe", x"03",
    x"f6", x"fd", x"00", x"f3", x"fe", x"03", x"ff", x"02",
    x"19", x"e6", x"02", x"c7", x"7f", x"46", x"c4", x"cc",
    x"09", x"39", x"c0", x"03", x"e3", x"fa", x"4d", x"1e",
    x"36", x"1c", x"1b", x"de", x"0f", x"15", x"b9", x"94",
    x"1e", x"f0", x"ec", x"35", x"60", x"12", x"fe", x"db",
    x"20", x"11", x"f1", x"2c", x"fe", x"e8", x"04", x"fd",
    x"28", x"fa", x"05", x"13", x"ab", x"da", x"ef", x"26",
    x"12", x"2a", x"15", x"05", x"c5", x"fa", x"e3", x"f6",
    x"07", x"f3", x"f3", x"d8", x"b2", x"dc", x"b9", x"ff",
    x"fa", x"06", x"01", x"02", x"fa", x"03", x"06", x"02",
    x"24", x"45", x"19", x"f5", x"fa", x"11", x"5a", x"16",
    x"0e", x"ff", x"01", x"02", x"fd", x"02", x"07", x"02",
    x"00", x"02", x"53", x"10", x"ef", x"0a", x"f5", x"28",
    x"cd", x"4b", x"3c", x"0a", x"07", x"f3", x"42", x"0b",
    x"13", x"0e", x"e9", x"eb", x"eb", x"e8", x"e0", x"df",
    x"9b", x"bf", x"3f", x"49", x"56", x"1d", x"0e", x"fc",
    x"1b", x"d2", x"29", x"1a", x"7a", x"45", x"d7", x"01",
    x"f5", x"c6", x"2a", x"f2", x"03", x"1e", x"41", x"fd",
    x"10", x"4d", x"a3", x"ca", x"da", x"e9", x"b1", x"d4",
    x"d4", x"ff", x"06", x"ef", x"11", x"25", x"0c", x"f9",
    x"f5", x"c9", x"0f", x"3a", x"0f", x"2c", x"c4", x"f5",
    x"b8", x"bf", x"aa", x"a9", x"16", x"37", x"e7", x"39",
    x"f6", x"ff", x"2d", x"f5", x"01", x"32", x"fb", x"2b",
    x"c5", x"cf", x"e2", x"d4", x"48", x"c9", x"4d", x"df",
    x"9b", x"25", x"f4", x"f4", x"1a", x"13", x"e8", x"f5",
    x"a3", x"1f", x"28", x"2e", x"11", x"fa", x"52", x"37",
    x"0d", x"e3", x"ba", x"05", x"35", x"50", x"41", x"1d",
    x"f0", x"f7", x"19", x"41", x"44", x"fe", x"2a", x"f6",
    x"02", x"1f", x"2b", x"41", x"0c", x"09", x"4f", x"32",
    x"2b", x"31", x"35", x"30", x"16", x"f9", x"09", x"bf",
    x"ed", x"02", x"00", x"01", x"23", x"05", x"07", x"e3",
    x"07", x"d3", x"1f", x"b3", x"fd", x"06", x"aa", x"07",
    x"ea", x"30", x"0c", x"d6", x"17", x"17", x"f6", x"cb",
    x"07", x"15", x"74", x"3f", x"fe", x"27", x"1f", x"23",
    x"e5", x"e3", x"1d", x"de", x"ed", x"21", x"e8", x"ae",
    x"b7", x"f7", x"6d", x"87", x"ec", x"c1", x"f3", x"58",
    x"9f", x"f0", x"9a", x"1c", x"08", x"e9", x"0e", x"1e",
    x"1f", x"f4", x"f5", x"3e", x"02", x"25", x"26", x"fa",
    x"d3", x"0d", x"ca", x"01", x"1d", x"fa", x"21", x"e2",
    x"4c", x"5e", x"e8", x"1b", x"32", x"eb", x"1b", x"3a",
    x"73", x"dd", x"36", x"f0", x"fc", x"08", x"29", x"f6",
    x"a6", x"0b", x"f3", x"51", x"29", x"ef", x"35", x"0a",
    x"ce", x"35", x"c7", x"1f", x"1b", x"ed", x"04", x"ea",
    x"f1", x"fc", x"ec", x"ea", x"bd", x"00", x"fc", x"d3",
    x"0e", x"21", x"f0", x"df", x"9a", x"d4", x"cc", x"06",
    x"06", x"04", x"00", x"01", x"fe", x"04", x"00", x"00",
    x"f8", x"fe", x"f2", x"0b", x"94", x"c2", x"15", x"ec",
    x"b6", x"01", x"07", x"00", x"fc", x"fc", x"00", x"f9",
    x"04", x"fb", x"22", x"17", x"11", x"b8", x"f0", x"f8",
    x"07", x"0a", x"00", x"08", x"00", x"d2", x"e5", x"f0",
    x"fa", x"f0", x"18", x"17", x"1e", x"0c", x"01", x"41",
    x"d1", x"2c", x"3f", x"99", x"3e", x"25", x"fe", x"1e",
    x"1c", x"ee", x"ff", x"0b", x"3c", x"51", x"15", x"46",
    x"a0", x"f8", x"55", x"d2", x"40", x"1a", x"0f", x"39",
    x"f2", x"11", x"2f", x"1f", x"df", x"27", x"e8", x"d3",
    x"f9", x"27", x"1c", x"35", x"35", x"0b", x"9d", x"0a",
    x"f4", x"3d", x"f5", x"3f", x"f2", x"d0", x"0b", x"20",
    x"e0", x"03", x"ef", x"e9", x"1a", x"03", x"2f", x"07",
    x"01", x"ea", x"15", x"19", x"fb", x"f3", x"20", x"f3",
    x"0f", x"08", x"af", x"de", x"da", x"ff", x"fb", x"06",
    x"c3", x"c2", x"c8", x"ab", x"0a", x"f1", x"ec", x"25",
    x"1c", x"e8", x"e5", x"ba", x"fb", x"26", x"38", x"0c",
    x"0f", x"f2", x"c6", x"14", x"57", x"94", x"0c", x"ec",
    x"f8", x"ff", x"e9", x"0f", x"2e", x"e8", x"f2", x"3d",
    x"21", x"cb", x"0d", x"01", x"08", x"26", x"a7", x"15",
    x"58", x"e4", x"e2", x"d0", x"0c", x"f4", x"d4", x"2a",
    x"cc", x"de", x"1f", x"01", x"2f", x"f2", x"e3", x"ff",
    x"b1", x"11", x"52", x"06", x"1b", x"17", x"f0", x"04",
    x"1c", x"e7", x"df", x"d8", x"fa", x"e4", x"02", x"fe",
    x"ca", x"35", x"bb", x"1a", x"3d", x"01", x"dc", x"f7",
    x"0e", x"22", x"14", x"34", x"f6", x"2f", x"25", x"e4",
    x"fa", x"da", x"b9", x"aa", x"bd", x"bb", x"e3", x"09",
    x"f6", x"25", x"08", x"0d", x"ec", x"11", x"e9", x"14",
    x"be", x"84", x"e8", x"33", x"10", x"11", x"14", x"e7",
    x"10", x"19", x"be", x"be", x"15", x"30", x"30", x"e0",
    x"ff", x"ad", x"dc", x"05", x"08", x"b8", x"04", x"17",
    x"32", x"23", x"fe", x"f1", x"da", x"b8", x"29", x"12",
    x"01", x"22", x"df", x"fc", x"bd", x"d2", x"07", x"e9",
    x"fa", x"24", x"b0", x"ea", x"00", x"d5", x"c2", x"cd",
    x"e7", x"11", x"2d", x"ed", x"f9", x"04", x"09", x"02",
    x"1f", x"4e", x"0f", x"44", x"cf", x"d0", x"ba", x"fc",
    x"07", x"05", x"ff", x"ff", x"fe", x"fd", x"fd", x"05",
    x"14", x"1a", x"e9", x"04", x"7e", x"bb", x"cd", x"ea",
    x"46", x"fc", x"fa", x"02", x"05", x"fd", x"fd", x"ff",
    x"fe", x"fa", x"f0", x"e9", x"c3", x"f2", x"b0", x"d9",
    x"ed", x"2a", x"f9", x"f4", x"ca", x"0c", x"d6", x"fa",
    x"1d", x"20", x"2c", x"e4", x"e2", x"06", x"04", x"2d",
    x"db", x"1e", x"1a", x"1e", x"00", x"0d", x"04", x"bf",
    x"0f", x"46", x"03", x"cd", x"e3", x"f9", x"0e", x"02",
    x"1b", x"51", x"00", x"2b", x"ad", x"d6", x"d5", x"dd",
    x"a3", x"b6", x"e8", x"17", x"fb", x"cb", x"ff", x"e9",
    x"aa", x"08", x"08", x"16", x"34", x"05", x"b7", x"04",
    x"fb", x"01", x"e4", x"b5", x"0d", x"06", x"08", x"03",
    x"21", x"41", x"94", x"94", x"94", x"1f", x"22", x"3f",
    x"25", x"2d", x"c7", x"75", x"13", x"fb", x"ed", x"37",
    x"19", x"cb", x"c2", x"f6", x"e8", x"f5", x"1c", x"e4",
    x"39", x"d4", x"f2", x"e5", x"d6", x"ec", x"03", x"05",
    x"0e", x"0b", x"05", x"5e", x"97", x"e4", x"c6", x"f7",
    x"2d", x"4b", x"0e", x"03", x"28", x"d6", x"04", x"0f",
    x"24", x"b2", x"b1", x"e2", x"b5", x"d5", x"e4", x"d9",
    x"f3", x"c3", x"fc", x"2b", x"1f", x"2e", x"1b", x"20",
    x"4c", x"0d", x"d6", x"e8", x"45", x"13", x"13", x"d9",
    x"92", x"8f", x"0f", x"eb", x"c4", x"19", x"ff", x"18",
    x"f8", x"f1", x"1f", x"a2", x"59", x"ea", x"15", x"09",
    x"21", x"11", x"fc", x"04", x"c7", x"88", x"dc", x"19",
    x"2f", x"29", x"d1", x"f5", x"0a", x"d6", x"96", x"af",
    x"14", x"10", x"4a", x"12", x"06", x"fb", x"f5", x"dc",
    x"f5", x"ec", x"d0", x"c0", x"e0", x"f2", x"01", x"ad",
    x"9a", x"d7", x"0b", x"14", x"fe", x"0d", x"12", x"c8",
    x"e0", x"c5", x"c3", x"b3", x"0a", x"22", x"ed", x"b2",
    x"0f", x"04", x"f2", x"2c", x"22", x"0e", x"37", x"1e",
    x"0b", x"45", x"07", x"30", x"1a", x"28", x"27", x"49",
    x"f3", x"03", x"3e", x"d3", x"15", x"16", x"1d", x"1d",
    x"0c", x"22", x"14", x"16", x"e2", x"9f", x"a5", x"ec",
    x"0e", x"fe", x"e0", x"fb", x"f6", x"e0", x"c2", x"e1",
    x"ed", x"eb", x"eb", x"06", x"1d", x"01", x"96", x"03",
    x"f7", x"f3", x"17", x"17", x"20", x"29", x"1b", x"ff",
    x"fe", x"fc", x"fc", x"01", x"fa", x"06", x"fb", x"07",
    x"1a", x"16", x"0b", x"05", x"e8", x"11", x"40", x"e5",
    x"11", x"fd", x"00", x"fd", x"fe", x"fc", x"fc", x"06",
    x"02", x"03", x"ef", x"f9", x"cb", x"1f", x"f8", x"da",
    x"0e", x"39", x"00", x"c5", x"ba", x"d3", x"de", x"0c",
    x"f9", x"f6", x"e1", x"bd", x"1a", x"f6", x"e1", x"50",
    x"0b", x"07", x"2e", x"28", x"1d", x"da", x"ec", x"05",
    x"0e", x"2d", x"1b", x"12", x"0b", x"f0", x"07", x"1c",
    x"b5", x"67", x"0b", x"0e", x"e0", x"20", x"1b", x"eb",
    x"28", x"23", x"ec", x"0e", x"19", x"e8", x"fa", x"0c",
    x"e4", x"d7", x"c2", x"15", x"17", x"21", x"2b", x"29",
    x"4b", x"1e", x"de", x"0d", x"21", x"11", x"f2", x"e5",
    x"11", x"31", x"e2", x"d9", x"cb", x"f8", x"02", x"10",
    x"13", x"08", x"18", x"05", x"e5", x"97", x"3d", x"f3",
    x"c2", x"2d", x"01", x"f7", x"fc", x"02", x"2b", x"f2",
    x"19", x"1f", x"51", x"38", x"f7", x"da", x"fe", x"f2",
    x"0b", x"2a", x"00", x"27", x"25", x"24", x"09", x"f0",
    x"ce", x"15", x"37", x"1b", x"1c", x"2a", x"0b", x"e5",
    x"c3", x"8e", x"11", x"2c", x"bc", x"0d", x"09", x"fd",
    x"50", x"37", x"18", x"54", x"13", x"06", x"0c", x"0a",
    x"1d", x"fd", x"02", x"9e", x"e7", x"f9", x"ee", x"1a",
    x"d7", x"07", x"fd", x"ff", x"ef", x"07", x"fb", x"f8",
    x"d7", x"07", x"4d", x"2e", x"21", x"c2", x"2d", x"ea",
    x"c3", x"fb", x"cd", x"ea", x"13", x"df", x"f7", x"ff",
    x"f2", x"de", x"1d", x"19", x"fb", x"f7", x"f0", x"f3",
    x"d3", x"f9", x"1f", x"c9", x"0a", x"19", x"2a", x"07",
    x"f4", x"e1", x"e1", x"d7", x"ce", x"d6", x"e4", x"ee",
    x"b7", x"ca", x"1c", x"d1", x"e0", x"02", x"e2", x"f5",
    x"f1", x"5b", x"42", x"d0", x"fa", x"dc", x"90", x"08",
    x"01", x"ab", x"2f", x"e5", x"94", x"16", x"e2", x"c7",
    x"ac", x"0d", x"03", x"f3", x"42", x"25", x"e2", x"07",
    x"10", x"d1", x"d0", x"0b", x"d5", x"d3", x"a6", x"d9",
    x"ce", x"b2", x"f0", x"fc", x"f0", x"31", x"fc", x"e8",
    x"d8", x"9f", x"14", x"3b", x"22", x"11", x"c8", x"eb",
    x"d7", x"db", x"ff", x"14", x"03", x"0b", x"94", x"c4",
    x"c0", x"f2", x"f2", x"f0", x"f2", x"e9", x"01", x"01",
    x"05", x"07", x"05", x"ff", x"01", x"fa", x"f9", x"05",
    x"e9", x"e3", x"0d", x"05", x"14", x"70", x"2f", x"21",
    x"d2", x"ff", x"fa", x"04", x"ff", x"02", x"06", x"03",
    x"05", x"fb", x"24", x"50", x"19", x"03", x"f3", x"de",
    x"3b", x"02", x"c2", x"11", x"2e", x"23", x"cd", x"cb",
    x"c9", x"cb", x"b8", x"ed", x"bf", x"12", x"de", x"ea",
    x"0e", x"08", x"de", x"0b", x"f0", x"f3", x"24", x"f3",
    x"c0", x"00", x"34", x"24", x"f3", x"ee", x"0c", x"e9",
    x"03", x"11", x"f8", x"e4", x"c2", x"00", x"c0", x"14",
    x"fe", x"2f", x"ff", x"50", x"32", x"8a", x"fc", x"fd",
    x"d6", x"b6", x"06", x"d2", x"00", x"0d", x"3b", x"f9",
    x"f3", x"25", x"04", x"dc", x"11", x"e3", x"e5", x"1e",
    x"0d", x"f4", x"fb", x"12", x"eb", x"55", x"9a", x"9d",
    x"75", x"f4", x"02", x"e9", x"ec", x"eb", x"d9", x"8f",
    x"d0", x"d1", x"fa", x"fb", x"aa", x"ad", x"f2", x"0a",
    x"f1", x"09", x"d0", x"0c", x"11", x"eb", x"f4", x"fc",
    x"c2", x"f2", x"f7", x"19", x"29", x"19", x"0d", x"2c",
    x"05", x"d4", x"f6", x"0d", x"a5", x"13", x"ef", x"09",
    x"09", x"03", x"ee", x"e3", x"c7", x"64", x"ca", x"be",
    x"2b", x"fc", x"f0", x"e9", x"fa", x"ea", x"cb", x"f0",
    x"e9", x"1c", x"0c", x"db", x"5e", x"85", x"a2", x"22",
    x"00", x"04", x"14", x"0f", x"bd", x"f2", x"0b", x"e8",
    x"4c", x"29", x"17", x"e2", x"ed", x"eb", x"c9", x"bb",
    x"88", x"06", x"36", x"fc", x"ec", x"0c", x"e4", x"a5",
    x"f6", x"dd", x"e8", x"21", x"db", x"31", x"33", x"24",
    x"e9", x"e4", x"74", x"8f", x"db", x"d9", x"fd", x"11",
    x"11", x"ec", x"12", x"f4", x"f8", x"e5", x"ef", x"0e",
    x"05", x"30", x"cc", x"e1", x"04", x"b7", x"18", x"02",
    x"11", x"f4", x"c9", x"07", x"e9", x"f4", x"15", x"09",
    x"1a", x"2c", x"2c", x"ef", x"0c", x"cc", x"e8", x"e9",
    x"d1", x"e4", x"f3", x"00", x"cd", x"20", x"f5", x"f6",
    x"d8", x"0a", x"36", x"e7", x"db", x"f8", x"17", x"1c",
    x"1d", x"4b", x"0e", x"0d", x"ce", x"fe", x"4b", x"16",
    x"3b", x"c6", x"19", x"f0", x"bc", x"da", x"f7", x"16",
    x"49", x"30", x"fa", x"02", x"19", x"11", x"ef", x"e7",
    x"d3", x"fa", x"c6", x"2b", x"dd", x"f5", x"4d", x"ff",
    x"fe", x"01", x"fb", x"fc", x"00", x"04", x"fd", x"fa",
    x"c5", x"dc", x"b6", x"c9", x"d1", x"fb", x"0b", x"13",
    x"ff", x"03", x"fe", x"ff", x"ff", x"fd", x"05", x"05",
    x"02", x"fa", x"17", x"f9", x"fc", x"1d", x"e5", x"89",
    x"e0", x"df", x"b1", x"2a", x"3a", x"f0", x"e3", x"db",
    x"8c", x"dc", x"ea", x"29", x"d5", x"d0", x"ef", x"0a",
    x"39", x"21", x"2f", x"0a", x"c1", x"6c", x"82", x"7d",
    x"1e", x"20", x"12", x"0d", x"0e", x"92", x"95", x"d9",
    x"26", x"d4", x"16", x"0e", x"12", x"02", x"33", x"2b",
    x"16", x"20", x"d3", x"77", x"1d", x"1f", x"0b", x"e5",
    x"e1", x"e3", x"de", x"2f", x"01", x"a1", x"e3", x"0c",
    x"31", x"d2", x"e6", x"e2", x"3c", x"0c", x"df", x"26",
    x"de", x"14", x"da", x"02", x"b7", x"1e", x"14", x"a0",
    x"02", x"13", x"f5", x"31", x"e4", x"15", x"d7", x"1f",
    x"f6", x"f1", x"10", x"d6", x"0d", x"19", x"d0", x"09",
    x"29", x"73", x"09", x"f3", x"2b", x"b4", x"e4", x"fb",
    x"35", x"ee", x"df", x"1a", x"a7", x"12", x"1a", x"ae",
    x"bd", x"ee", x"14", x"fe", x"f6", x"f5", x"68", x"9e",
    x"b3", x"25", x"d3", x"00", x"c1", x"fd", x"04", x"ef",
    x"c4", x"2f", x"86", x"1d", x"25", x"78", x"46", x"ef",
    x"94", x"d7", x"d8", x"94", x"db", x"d7", x"a3", x"ce",
    x"cb", x"0d", x"a1", x"d7", x"f2", x"42", x"ef", x"66",
    x"30", x"9b", x"bf", x"f8", x"fc", x"1c", x"23", x"f6",
    x"ed", x"fd", x"ea", x"e2", x"d9", x"05", x"fb", x"35",
    x"1e", x"22", x"1b", x"f8", x"d4", x"0d", x"24", x"cd",
    x"36", x"f6", x"d9", x"d9", x"b0", x"a2", x"b3", x"e1",
    x"a9", x"17", x"ed", x"e4", x"f5", x"d1", x"d5", x"fc",
    x"b9", x"1c", x"05", x"02", x"1f", x"04", x"14", x"de",
    x"cc", x"b3", x"b7", x"f5", x"c0", x"c4", x"ff", x"dd",
    x"80", x"0b", x"7d", x"fa", x"63", x"70", x"3c", x"31",
    x"b5", x"d3", x"50", x"9f", x"ff", x"42", x"ed", x"2f",
    x"2e", x"34", x"25", x"e7", x"bd", x"e4", x"e8", x"c3",
    x"ce", x"16", x"d9", x"cf", x"06", x"d3", x"70", x"09",
    x"b5", x"fe", x"dc", x"91", x"02", x"0b", x"06", x"ab",
    x"d2", x"d8", x"2f", x"98", x"dd", x"18", x"ed", x"12",
    x"01", x"ba", x"f4", x"1c", x"be", x"13", x"d7", x"ff",
    x"07", x"fe", x"fe", x"fc", x"02", x"02", x"01", x"02",
    x"16", x"b4", x"9d", x"0b", x"a2", x"2e", x"0e", x"e8",
    x"fd", x"fe", x"02", x"fd", x"f9", x"00", x"f9", x"06",
    x"01", x"05", x"06", x"e0", x"59", x"1c", x"2b", x"11",
    x"1d", x"27", x"c3", x"05", x"74", x"a7", x"07", x"a3",
    x"0e", x"2d", x"ab", x"e8", x"3d", x"0e", x"f0", x"11",
    x"fa", x"1e", x"ff", x"fb", x"1b", x"d4", x"72", x"fa",
    x"20", x"bf", x"09", x"1e", x"1d", x"f3", x"1f", x"1a",
    x"ca", x"e0", x"21", x"b7", x"dd", x"f6", x"04", x"bd",
    x"f0", x"c4", x"e6", x"d2", x"b5", x"f0", x"07", x"e9",
    x"1b", x"ea", x"ca", x"c0", x"97", x"27", x"f2", x"0d",
    x"07", x"0f", x"fa", x"ac", x"eb", x"a5", x"06", x"dd",
    x"14", x"47", x"f7", x"2d", x"ec", x"f1", x"c7", x"09",
    x"ba", x"b7", x"ea", x"25", x"aa", x"b7", x"0b", x"2d",
    x"81", x"f1", x"da", x"eb", x"1b", x"17", x"07", x"4e",
    x"ed", x"cd", x"30", x"0c", x"89", x"fd", x"00", x"f5",
    x"ee", x"02", x"0a", x"07", x"a6", x"f1", x"4b", x"13",
    x"a9", x"3b", x"21", x"ab", x"21", x"f9", x"96", x"e9",
    x"3a", x"0f", x"09", x"c7", x"1d", x"37", x"50", x"16",
    x"14", x"1e", x"e3", x"0a", x"c9", x"15", x"18", x"a9",
    x"16", x"ba", x"07", x"92", x"d6", x"b4", x"23", x"f8",
    x"95", x"17", x"06", x"e1", x"bd", x"fb", x"e9", x"1f",
    x"1f", x"e1", x"de", x"f3", x"b0", x"f7", x"f7", x"c0",
    x"af", x"a8", x"9e", x"0f", x"21", x"d5", x"e2", x"e4",
    x"f8", x"07", x"d4", x"22", x"19", x"ca", x"b2", x"68",
    x"e5", x"83", x"87", x"11", x"b5", x"45", x"04", x"fa",
    x"fd", x"fa", x"f9", x"03", x"07", x"f5", x"fc", x"fc",
    x"85", x"ad", x"08", x"1c", x"a3", x"cc", x"ef", x"d7",
    x"ef", x"ff", x"f0", x"a1", x"f7", x"02", x"9a", x"0d",
    x"99", x"f9", x"22", x"0e", x"f9", x"07", x"44", x"e7",
    x"fe", x"47", x"16", x"52", x"15", x"e5", x"e1", x"14",
    x"68", x"1d", x"31", x"14", x"03", x"39", x"05", x"f6",
    x"ca", x"f9", x"ca", x"cf", x"13", x"01", x"f5", x"1b",
    x"f1", x"00", x"08", x"2b", x"fa", x"f9", x"3f", x"33",
    x"fe", x"ee", x"01", x"0c", x"bc", x"e9", x"1b", x"ca",
    x"d2", x"03", x"c2", x"ea", x"1c", x"13", x"ee", x"05",
    x"f9", x"f9", x"fa", x"fe", x"fe", x"fb", x"01", x"fc",
    x"ed", x"db", x"e9", x"db", x"e7", x"e4", x"89", x"12",
    x"1a", x"fb", x"06", x"04", x"01", x"00", x"06", x"05",
    x"04", x"fa", x"08", x"13", x"18", x"f9", x"1c", x"ea",
    x"17", x"49", x"27", x"25", x"13", x"50", x"f0", x"8d",
    x"0c", x"f7", x"f4", x"3f", x"33", x"48", x"23", x"eb",
    x"b4", x"c5", x"40", x"39", x"d5", x"1b", x"f2", x"dd",
    x"e3", x"d3", x"e8", x"1e", x"30", x"df", x"08", x"2e",
    x"10", x"e7", x"19", x"d1", x"f5", x"26", x"fc", x"29",
    x"3e", x"28", x"e3", x"15", x"f1", x"b7", x"cd", x"82",
    x"10", x"26", x"2c", x"ee", x"14", x"49", x"02", x"cc",
    x"10", x"fb", x"1b", x"22", x"e0", x"ce", x"00", x"00",
    x"07", x"fe", x"d8", x"05", x"0d", x"03", x"d7", x"0d",
    x"0c", x"86", x"ea", x"0a", x"06", x"31", x"10", x"ee",
    x"cb", x"12", x"27", x"f3", x"1a", x"02", x"1b", x"fd",
    x"ed", x"2e", x"dc", x"11", x"f7", x"bc", x"73", x"da",
    x"fa", x"37", x"fa", x"59", x"61", x"ee", x"10", x"0b",
    x"e6", x"12", x"29", x"e5", x"3f", x"3b", x"43", x"e4",
    x"e6", x"17", x"27", x"25", x"1e", x"f7", x"04", x"f5",
    x"e9", x"00", x"ed", x"ec", x"e8", x"d6", x"15", x"1b",
    x"fd", x"ff", x"f1", x"db", x"f9", x"d2", x"b8", x"dc",
    x"c2", x"e6", x"0f", x"02", x"fa", x"da", x"e9", x"0b",
    x"27", x"14", x"21", x"f2", x"d8", x"e6", x"f7", x"f5",
    x"09", x"fc", x"dc", x"9e", x"3f", x"19", x"1f", x"32",
    x"26", x"3b", x"02", x"22", x"fb", x"f4", x"1f", x"4f",
    x"c6", x"d1", x"27", x"e5", x"fd", x"27", x"f9", x"f4",
    x"f6", x"d6", x"d4", x"c8", x"07", x"fe", x"e5", x"fc",
    x"29", x"16", x"ae", x"bf", x"06", x"09", x"12", x"c7",
    x"04", x"9c", x"1f", x"a5", x"a7", x"f7", x"eb", x"e2",
    x"dd", x"dd", x"2d", x"41", x"ca", x"0c", x"30", x"1b",
    x"e2", x"b0", x"0e", x"e3", x"18", x"e6", x"12", x"20",
    x"fa", x"01", x"ba", x"f7", x"f2", x"f4", x"37", x"f2",
    x"16", x"26", x"2e", x"08", x"f3", x"0a", x"db", x"0a",
    x"ef", x"14", x"fa", x"eb", x"00", x"e2", x"cb", x"eb",
    x"f0", x"f6", x"f8", x"d9", x"3d", x"07", x"f3", x"9e",
    x"cf", x"d5", x"fa", x"f6", x"18", x"f5", x"b0", x"02",
    x"04", x"03", x"04", x"fb", x"fc", x"fe", x"05", x"06",
    x"11", x"da", x"f2", x"ea", x"9c", x"ad", x"f5", x"c8",
    x"de", x"fe", x"f9", x"05", x"fd", x"ff", x"fb", x"03",
    x"fa", x"fc", x"16", x"3f", x"0d", x"ed", x"23", x"eb",
    x"cc", x"0f", x"b8", x"08", x"d1", x"d0", x"02", x"55",
    x"46", x"20", x"f0", x"a6", x"2a", x"03", x"57", x"2a",
    x"11", x"4a", x"4c", x"2c", x"41", x"f7", x"04", x"1e",
    x"0b", x"12", x"ee", x"0f", x"fd", x"11", x"42", x"2a",
    x"ee", x"ff", x"f8", x"dd", x"3a", x"25", x"14", x"fe",
    x"e5", x"21", x"33", x"05", x"53", x"da", x"1d", x"4b",
    x"eb", x"fa", x"1d", x"0b", x"1a", x"d7", x"10", x"17",
    x"66", x"f3", x"0f", x"3d", x"09", x"d6", x"01", x"f4",
    x"1f", x"e0", x"fc", x"8f", x"d6", x"cb", x"a2", x"05",
    x"07", x"25", x"23", x"f0", x"ff", x"15", x"d3", x"26",
    x"ab", x"5b", x"30", x"e1", x"d8", x"79", x"ed", x"03",
    x"e4", x"e7", x"f2", x"21", x"9a", x"08", x"04", x"26",
    x"d7", x"11", x"24", x"18", x"0b", x"f6", x"1a", x"13",
    x"09", x"05", x"04", x"0c", x"21", x"dc", x"10", x"25",
    x"ec", x"14", x"29", x"07", x"1f", x"1f", x"e6", x"f5",
    x"05", x"14", x"3b", x"13", x"34", x"3f", x"f7", x"2a",
    x"4f", x"d3", x"7d", x"bd", x"e9", x"b0", x"fd", x"3a",
    x"12", x"74", x"04", x"d1", x"2a", x"18", x"e4", x"35",
    x"fc", x"c9", x"1d", x"1d", x"dd", x"fb", x"dd", x"00",
    x"00", x"18", x"07", x"cd", x"0e", x"0a", x"57", x"17",
    x"f5", x"20", x"f3", x"04", x"32", x"de", x"f6", x"6b",
    x"cc", x"ea", x"17", x"00", x"d2", x"d2", x"e9", x"cf",
    x"14", x"ed", x"f8", x"f9", x"c8", x"ca", x"ca", x"dd",
    x"a8", x"ef", x"c0", x"f0", x"c8", x"14", x"10", x"04",
    x"d4", x"df", x"dc", x"f1", x"f0", x"e1", x"0b", x"0d",
    x"28", x"37", x"2f", x"f4", x"d8", x"d0", x"07", x"d3",
    x"25", x"26", x"d9", x"07", x"3b", x"09", x"00", x"fe",
    x"f4", x"d6", x"02", x"06", x"f7", x"bd", x"ea", x"f8",
    x"f3", x"1d", x"eb", x"fb", x"db", x"e8", x"f8", x"05",
    x"05", x"e6", x"31", x"19", x"35", x"d0", x"04", x"f2",
    x"f9", x"18", x"1e", x"18", x"06", x"fb", x"2f", x"bf",
    x"f1", x"09", x"18", x"fe", x"10", x"2e", x"00", x"f9",
    x"06", x"02", x"05", x"fb", x"fc", x"fb", x"05", x"04",
    x"4d", x"f8", x"0b", x"12", x"04", x"21", x"0b", x"cc",
    x"f8", x"f9", x"fe", x"fe", x"f9", x"03", x"fb", x"07",
    x"00", x"fd", x"fb", x"16", x"ab", x"da", x"09", x"fd",
    x"03", x"b4", x"e2", x"f5", x"f3", x"ed", x"1b", x"d7",
    x"90", x"05", x"1d", x"e1", x"fb", x"f6", x"1f", x"09",
    x"d0", x"12", x"2b", x"b1", x"fd", x"3f", x"20", x"0a",
    x"e6", x"c1", x"09", x"f1", x"0d", x"31", x"20", x"27",
    x"04", x"16", x"05", x"ee", x"1a", x"29", x"0a", x"82",
    x"fa", x"05", x"15", x"33", x"05", x"68", x"c0", x"da",
    x"e4", x"20", x"3d", x"e9", x"fb", x"fe", x"d4", x"20",
    x"29", x"fe", x"00", x"2f", x"09", x"e4", x"0b", x"04",
    x"ef", x"15", x"d2", x"f1", x"d0", x"64", x"d6", x"24",
    x"4d", x"03", x"52", x"c2", x"e9", x"e8", x"f6", x"0a",
    x"e5", x"41", x"05", x"f3", x"fc", x"f7", x"f7", x"04",
    x"00", x"31", x"0c", x"03", x"f8", x"fb", x"f2", x"18",
    x"31", x"06", x"01", x"31", x"f4", x"1f", x"e3", x"04",
    x"2f", x"dd", x"ff", x"15", x"1a", x"08", x"1e", x"f3",
    x"18", x"1a", x"ec", x"0e", x"40", x"fc", x"f9", x"f2",
    x"db", x"f1", x"4b", x"00", x"18", x"3c", x"3f", x"4e",
    x"01", x"24", x"b7", x"af", x"10", x"03", x"c7", x"e2",
    x"0c", x"56", x"ed", x"28", x"1c", x"cf", x"b4", x"00",
    x"d5", x"e9", x"15", x"ea", x"e2", x"dd", x"f7", x"fb",
    x"68", x"31", x"42", x"45", x"bd", x"f4", x"23", x"f3",
    x"2c", x"2a", x"1d", x"38", x"0d", x"25", x"1d", x"c9",
    x"f2", x"dc", x"db", x"1c", x"ce", x"ca", x"fc", x"dc",
    x"f5", x"e7", x"fd", x"f0", x"a5", x"a4", x"5c", x"e8",
    x"00", x"dd", x"20", x"d3", x"d8", x"50", x"0b", x"17",
    x"f9", x"1f", x"1d", x"ea", x"35", x"36", x"28", x"2b",
    x"24", x"22", x"3f", x"4d", x"fe", x"ed", x"db", x"fb",
    x"db", x"2c", x"ce", x"b4", x"08", x"e2", x"d0", x"e5",
    x"9f", x"c3", x"c9", x"20", x"db", x"06", x"2c", x"ef",
    x"2f", x"b0", x"c2", x"f4", x"fe", x"12", x"21", x"f7",
    x"0b", x"1d", x"d5", x"ea", x"8d", x"eb", x"07", x"0d",
    x"00", x"0c", x"21", x"90", x"c4", x"d1", x"16", x"fc",
    x"d6", x"22", x"eb", x"a3", x"21", x"35", x"ee", x"fb",
    x"00", x"fb", x"05", x"07", x"06", x"f9", x"03", x"ff",
    x"18", x"1b", x"f0", x"ec", x"de", x"f9", x"05", x"14",
    x"dd", x"fc", x"fc", x"05", x"fc", x"fe", x"fc", x"04",
    x"fd", x"fc", x"08", x"0c", x"44", x"31", x"fd", x"03",
    x"24", x"ed", x"ea", x"0a", x"ec", x"15", x"1a", x"da",
    x"97", x"16", x"e6", x"db", x"f5", x"a8", x"f3", x"3f",
    x"57", x"27", x"9d", x"e7", x"cc", x"25", x"f4", x"41",
    x"31", x"12", x"f5", x"fa", x"d9", x"12", x"16", x"08",
    x"e2", x"13", x"d2", x"20", x"fa", x"e0", x"d5", x"e9",
    x"da", x"cb", x"24", x"f4", x"33", x"df", x"08", x"2e",
    x"e3", x"28", x"11", x"12", x"e9", x"f1", x"b9", x"e2",
    x"05", x"07", x"19", x"08", x"ec", x"e1", x"cb", x"48",
    x"80", x"4f", x"d4", x"b9", x"0a", x"1d", x"22", x"08",
    x"1f", x"24", x"c8", x"db", x"18", x"12", x"40", x"22",
    x"1e", x"e1", x"cd", x"84", x"d6", x"e2", x"cc", x"1a",
    x"f7", x"c7", x"ef", x"b4", x"d7", x"06", x"10", x"14",
    x"25", x"1f", x"05", x"3f", x"00", x"e5", x"dd", x"00",
    x"ea", x"0f", x"f7", x"e1", x"47", x"f8", x"f8", x"f9",
    x"f2", x"d7", x"37", x"f0", x"09", x"1b", x"1a", x"9a",
    x"df", x"f5", x"0b", x"f8", x"35", x"53", x"15", x"a2",
    x"77", x"fa", x"f5", x"10", x"3c", x"1c", x"05", x"37",
    x"0c", x"ed", x"2f", x"0d", x"15", x"f4", x"eb", x"c2",
    x"c3", x"64", x"13", x"ef", x"f6", x"ea", x"3d", x"10",
    x"1f", x"1f", x"1e", x"9d", x"d5", x"e3", x"03", x"28",
    x"15", x"3a", x"d7", x"db", x"30", x"fd", x"f0", x"0f",
    x"27", x"fc", x"f9", x"15", x"f0", x"b3", x"e4", x"93",
    x"b5", x"d9", x"8c", x"d9", x"e0", x"b0", x"de", x"fe",
    x"0e", x"d8", x"fb", x"08", x"19", x"1d", x"1d", x"09",
    x"1f", x"01", x"d0", x"16", x"05", x"d4", x"da", x"dd",
    x"21", x"09", x"f5", x"c4", x"1d", x"dc", x"1e", x"0e",
    x"06", x"d7", x"95", x"c8", x"e3", x"fc", x"19", x"2e",
    x"0b", x"03", x"16", x"07", x"32", x"de", x"03", x"07",
    x"0c", x"3d", x"20", x"38", x"24", x"ea", x"20", x"f6",
    x"ef", x"1d", x"d5", x"be", x"87", x"f9", x"2b", x"b6",
    x"c9", x"da", x"d3", x"4b", x"0d", x"f2", x"f7", x"d0",
    x"ef", x"fb", x"ef", x"f4", x"01", x"df", x"c4", x"fb",
    x"fa", x"ff", x"ff", x"f9", x"05", x"06", x"fd", x"fd",
    x"18", x"0a", x"37", x"e7", x"cb", x"da", x"f3", x"18",
    x"c5", x"02", x"f9", x"03", x"fe", x"fd", x"01", x"04",
    x"04", x"07", x"d7", x"bf", x"08", x"11", x"25", x"05",
    x"0d", x"18", x"33", x"f0", x"00", x"df", x"20", x"0c",
    x"1c", x"e5", x"c2", x"b1", x"2e", x"fe", x"e0", x"f6",
    x"07", x"3a", x"27", x"33", x"0c", x"09", x"3a", x"14",
    x"01", x"0b", x"1d", x"25", x"34", x"14", x"0d", x"f6",
    x"fa", x"c6", x"bd", x"e8", x"28", x"fe", x"ce", x"4a",
    x"0a", x"ff", x"e8", x"c8", x"e9", x"22", x"30", x"22",
    x"ff", x"b0", x"a2", x"ee", x"f4", x"e5", x"03", x"13",
    x"e1", x"0f", x"d6", x"ab", x"dd", x"00", x"1b", x"04",
    x"b2", x"fc", x"e5", x"ed", x"d4", x"b3", x"d0", x"49",
    x"37", x"5b", x"21", x"ee", x"da", x"f1", x"be", x"03",
    x"e6", x"de", x"cc", x"1f", x"15", x"2b", x"35", x"f6",
    x"ef", x"20", x"1a", x"0f", x"c8", x"0f", x"e9", x"1d",
    x"bc", x"f5", x"3b", x"1c", x"12", x"dd", x"05", x"fd",
    x"f1", x"e9", x"e2", x"e4", x"cc", x"0e", x"1c", x"2c",
    x"3f", x"17", x"17", x"ea", x"b4", x"fe", x"cf", x"ed",
    x"fc", x"ad", x"0a", x"f1", x"1e", x"52", x"3e", x"3b",
    x"5c", x"e5", x"fc", x"21", x"09", x"e9", x"d3", x"fa",
    x"f4", x"eb", x"15", x"f8", x"fd", x"b4", x"0b", x"1a",
    x"08", x"f3", x"a1", x"13", x"3b", x"13", x"21", x"a1",
    x"b3", x"bd", x"a0", x"77", x"20", x"2b", x"23", x"c3",
    x"de", x"fe", x"17", x"0c", x"0b", x"fb", x"c0", x"bf",
    x"16", x"e4", x"37", x"da", x"26", x"1b", x"d6", x"00",
    x"10", x"c2", x"f4", x"19", x"e5", x"f3", x"f8", x"03",
    x"0c", x"e8", x"fe", x"bf", x"c4", x"1e", x"29", x"f6",
    x"04", x"08", x"f3", x"d3", x"f6", x"0d", x"0c", x"22",
    x"1d", x"03", x"26", x"18", x"05", x"45", x"fe", x"27",
    x"ff", x"3b", x"ec", x"1d", x"25", x"f1", x"e6", x"98",
    x"e0", x"f3", x"fa", x"1e", x"38", x"33", x"11", x"18",
    x"33", x"24", x"f4", x"19", x"00", x"1e", x"e0", x"44",
    x"15", x"5d", x"ed", x"fe", x"ae", x"c4", x"ea", x"08",
    x"db", x"11", x"1c", x"f6", x"e4", x"3e", x"21", x"1f",
    x"01", x"a8", x"c6", x"10", x"c1", x"01", x"08", x"02",
    x"fd", x"fa", x"fc", x"01", x"03", x"06", x"ff", x"fe",
    x"e1", x"02", x"f3", x"13", x"10", x"04", x"11", x"0c",
    x"12", x"03", x"01", x"f9", x"03", x"05", x"00", x"fc",
    x"fd", x"fc", x"ee", x"31", x"0f", x"0f", x"0e", x"d7",
    x"bc", x"e4", x"db", x"fa", x"f0", x"f2", x"0c", x"e9",
    x"bb", x"0a", x"28", x"fd", x"be", x"3d", x"13", x"f0",
    x"35", x"2a", x"fa", x"fc", x"e4", x"1b", x"20", x"fa",
    x"32", x"02", x"9e", x"20", x"14", x"f4", x"ce", x"f5",
    x"de", x"d1", x"ff", x"0a", x"25", x"e8", x"06", x"b0",
    x"38", x"3b", x"93", x"0a", x"3a", x"e4", x"99", x"f4",
    x"eb", x"e2", x"05", x"e7", x"c2", x"69", x"0d", x"0a",
    x"0f", x"be", x"12", x"fe", x"08", x"e8", x"b7", x"ea",
    x"a3", x"90", x"24", x"25", x"0c", x"1c", x"04", x"2e",
    x"17", x"29", x"1a", x"0e", x"04", x"d8", x"10", x"1d",
    x"ff", x"23", x"2a", x"ed", x"fd", x"14", x"10", x"ee",
    x"2b", x"19", x"0e", x"15", x"0f", x"0c", x"05", x"00",
    x"43", x"f6", x"0c", x"3a", x"32", x"30", x"9f", x"fc",
    x"ee", x"10", x"40", x"d7", x"20", x"15", x"e3", x"de",
    x"a5", x"c1", x"f7", x"f5", x"bd", x"09", x"11", x"07",
    x"04", x"2c", x"0d", x"13", x"10", x"f3", x"04", x"3f",
    x"52", x"0f", x"23", x"c9", x"ec", x"25", x"17", x"03",
    x"4a", x"12", x"f0", x"24", x"aa", x"fb", x"f4", x"2b",
    x"0e", x"c0", x"c4", x"12", x"f1", x"d9", x"f4", x"0b",
    x"c9", x"39", x"0c", x"d8", x"b6", x"07", x"00", x"46",
    x"42", x"1d", x"06", x"cf", x"af", x"f2", x"e7", x"23",
    x"2a", x"fd", x"16", x"37", x"28", x"42", x"d8", x"e4",
    x"e1", x"b9", x"c3", x"cb", x"92", x"be", x"f1", x"fd",
    x"2f", x"1c", x"12", x"0f", x"09", x"31", x"e0", x"ed",
    x"03", x"c4", x"1c", x"e3", x"99", x"fb", x"f1", x"08",
    x"0d", x"9b", x"d7", x"4c", x"d7", x"e6", x"16", x"ba",
    x"a5", x"2f", x"83", x"18", x"12", x"db", x"f1", x"08",
    x"c4", x"4f", x"e6", x"2a", x"df", x"5e", x"16", x"f8",
    x"2f", x"02", x"d4", x"00", x"14", x"95", x"a6", x"0c",
    x"c7", x"f3", x"fe", x"40", x"ea", x"18", x"0d", x"33",
    x"12", x"1b", x"18", x"17", x"ef", x"d3", x"e2", x"e0",
    x"05", x"e0", x"ce", x"01", x"0e", x"e6", x"43", x"07",
    x"ff", x"fc", x"00", x"fa", x"f9", x"fc", x"06", x"01",
    x"33", x"ca", x"1f", x"06", x"0a", x"07", x"1d", x"21",
    x"1d", x"ff", x"07", x"06", x"02", x"fa", x"fa", x"02",
    x"00", x"f9", x"eb", x"55", x"e7", x"c1", x"d3", x"ed",
    x"17", x"11", x"20", x"04", x"a8", x"a0", x"c2", x"99",
    x"c6", x"04", x"c0", x"15", x"dd", x"11", x"5b", x"21",
    x"2d", x"29", x"36", x"25", x"06", x"bc", x"f7", x"0e",
    x"24", x"08", x"05", x"a7", x"e2", x"e8", x"ff", x"f8",
    x"0d", x"23", x"21", x"30", x"15", x"00", x"0b", x"ee",
    x"e7", x"70", x"fb", x"0c", x"53", x"a2", x"18", x"f8",
    x"a7", x"21", x"26", x"25", x"2c", x"eb", x"1f", x"cc",
    x"f8", x"c0", x"01", x"2a", x"e6", x"31", x"dc", x"ff",
    x"32", x"e6", x"36", x"b6", x"12", x"04", x"18", x"0a",
    x"e6", x"db", x"14", x"02", x"1d", x"42", x"0d", x"02",
    x"0f", x"24", x"26", x"2a", x"dd", x"07", x"16", x"0d",
    x"10", x"eb", x"13", x"2a", x"31", x"0c", x"1c", x"15",
    x"18", x"e7", x"df", x"fa", x"45", x"23", x"e8", x"e5",
    x"dd", x"50", x"ec", x"e7", x"1b", x"26", x"20", x"cf",
    x"b7", x"dd", x"94", x"0d", x"1b", x"d5", x"27", x"1e",
    x"d1", x"20", x"79", x"1c", x"26", x"3a", x"de", x"1f",
    x"26", x"d6", x"fd", x"e7", x"d2", x"e6", x"bf", x"10",
    x"fd", x"1f", x"8c", x"df", x"0e", x"cb", x"d4", x"ff",
    x"ce", x"f3", x"e6", x"ba", x"01", x"ff", x"c3", x"21",
    x"13", x"15", x"1f", x"21", x"dc", x"ff", x"38", x"07",
    x"22", x"0a", x"29", x"1e", x"06", x"ed", x"d2", x"40",
    x"ac", x"c0", x"ea", x"6e", x"c3", x"ec", x"de", x"01",
    x"02", x"f3", x"03", x"d9", x"ba", x"e8", x"bf", x"d8",
    x"be", x"0a", x"e2", x"cd", x"04", x"df", x"12", x"0d"
  );

  type conv2_bias_64_t is array (0 to 63) of std_logic_vector(7 downto 0);
  constant conv2_bias : conv2_bias_64_t := (
    x"06", x"ca", x"b9", x"13", x"bf", x"e3", x"e4", x"c8",
    x"dc", x"c3", x"fe", x"e4", x"b3", x"d0", x"9b", x"bf",
    x"cc", x"f8", x"e1", x"da", x"d8", x"c2", x"e3", x"c7",
    x"ec", x"f5", x"e5", x"f6", x"bb", x"e6", x"a2", x"b4",
    x"df", x"f6", x"cd", x"ee", x"f4", x"9d", x"dc", x"d9",
    x"f6", x"b7", x"d4", x"c0", x"c0", x"af", x"fe", x"e9",
    x"f9", x"f8", x"9f", x"b8", x"e8", x"b0", x"f8", x"db",
    x"ff", x"b6", x"c3", x"ae", x"e3", x"d4", x"ba", x"b3"
  );

  type conv2_activation_post_process_eps_1_t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant conv2_activation_post_process_eps : conv2_activation_post_process_eps_1_t := (
    x"00"
  );

  type conv2_activation_post_process_min_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant conv2_activation_post_process_min_val : conv2_activation_post_process_min_val__t := (
    x"1e"
  );

  type conv2_activation_post_process_max_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant conv2_activation_post_process_max_val : conv2_activation_post_process_max_val__t := (
    x"39"
  );

  type fc1_weight_128_576_t is array (0 to 73727) of std_logic_vector(7 downto 0);
  constant fc1_weight : fc1_weight_128_576_t := (
    x"0f", x"2a", x"f5", x"fa", x"25", x"24", x"f8", x"0d",
    x"70", x"00", x"00", x"16", x"0f", x"e9", x"1e", x"aa",
    x"f5", x"16", x"f4", x"fc", x"da", x"e7", x"03", x"d4",
    x"21", x"2a", x"d3", x"f3", x"f5", x"e7", x"f7", x"f8",
    x"eb", x"0e", x"1e", x"d4", x"ca", x"2d", x"12", x"0c",
    x"17", x"46", x"0a", x"4b", x"13", x"bc", x"ef", x"1d",
    x"a9", x"dd", x"f1", x"dd", x"ef", x"bd", x"1f", x"2e",
    x"0c", x"09", x"17", x"e6", x"eb", x"dd", x"db", x"16",
    x"03", x"36", x"e7", x"de", x"f8", x"e5", x"ee", x"1e",
    x"11", x"18", x"18", x"19", x"0b", x"21", x"12", x"0c",
    x"26", x"d6", x"14", x"1d", x"25", x"0c", x"e7", x"01",
    x"c7", x"f0", x"30", x"57", x"f5", x"f1", x"25", x"23",
    x"27", x"16", x"ef", x"fe", x"f1", x"00", x"01", x"1c",
    x"eb", x"d3", x"43", x"0e", x"63", x"0f", x"49", x"25",
    x"17", x"24", x"31", x"42", x"21", x"3d", x"ee", x"b2",
    x"20", x"ed", x"bb", x"2e", x"12", x"e8", x"39", x"10",
    x"de", x"06", x"f2", x"db", x"00", x"ff", x"d6", x"3b",
    x"fd", x"eb", x"fe", x"34", x"04", x"24", x"ed", x"00",
    x"1c", x"49", x"5e", x"02", x"1e", x"3f", x"d2", x"0a",
    x"3f", x"fb", x"05", x"fe", x"fb", x"ff", x"fc", x"05",
    x"05", x"fe", x"18", x"d6", x"19", x"66", x"70", x"7a",
    x"98", x"c6", x"fc", x"e0", x"d0", x"1a", x"fa", x"ca",
    x"1c", x"be", x"d2", x"0a", x"ee", x"f5", x"1a", x"fb",
    x"0c", x"b6", x"08", x"1e", x"25", x"f4", x"c3", x"ed",
    x"f1", x"09", x"12", x"ae", x"c4", x"ef", x"09", x"25",
    x"1d", x"e9", x"f7", x"15", x"c8", x"12", x"31", x"18",
    x"3d", x"1e", x"08", x"38", x"11", x"3c", x"71", x"35",
    x"46", x"62", x"37", x"d5", x"f7", x"0c", x"ea", x"12",
    x"06", x"c9", x"c9", x"d8", x"00", x"0b", x"1a", x"fc",
    x"ec", x"1a", x"dd", x"ed", x"02", x"e2", x"1d", x"27",
    x"c4", x"fe", x"06", x"fd", x"02", x"f9", x"fb", x"fd",
    x"00", x"fa", x"02", x"f7", x"0f", x"df", x"da", x"e1",
    x"da", x"0a", x"25", x"e8", x"0a", x"31", x"54", x"33",
    x"0a", x"0f", x"0c", x"fb", x"c3", x"f5", x"e8", x"a5",
    x"ed", x"02", x"c8", x"f5", x"f4", x"99", x"be", x"da",
    x"eb", x"11", x"24", x"22", x"08", x"e6", x"e7", x"f3",
    x"fa", x"45", x"1b", x"17", x"27", x"1a", x"22", x"25",
    x"08", x"24", x"e1", x"e4", x"03", x"f9", x"1e", x"10",
    x"e0", x"28", x"f8", x"1c", x"13", x"e2", x"f6", x"fe",
    x"c9", x"06", x"0f", x"3b", x"23", x"f9", x"b7", x"11",
    x"f3", x"f3", x"21", x"19", x"fe", x"f9", x"fc", x"00",
    x"f7", x"fd", x"ff", x"fb", x"fd", x"21", x"d5", x"df",
    x"f9", x"eb", x"f7", x"25", x"da", x"e2", x"09", x"47",
    x"04", x"e1", x"f2", x"ee", x"6d", x"d6", x"e7", x"13",
    x"25", x"f8", x"25", x"1c", x"15", x"0b", x"be", x"ba",
    x"fe", x"01", x"03", x"fb", x"00", x"fc", x"01", x"ff",
    x"04", x"0c", x"af", x"cb", x"8d", x"df", x"f8", x"0f",
    x"d7", x"fe", x"05", x"46", x"16", x"2a", x"16", x"26",
    x"93", x"d9", x"26", x"11", x"04", x"f2", x"a7", x"dd",
    x"17", x"53", x"37", x"33", x"b6", x"d3", x"c6", x"af",
    x"d7", x"f3", x"bc", x"da", x"f2", x"d9", x"53", x"70",
    x"1a", x"15", x"28", x"e8", x"14", x"0a", x"b1", x"33",
    x"4b", x"8b", x"db", x"24", x"d0", x"d2", x"0a", x"e6",
    x"86", x"09", x"e8", x"e5", x"dd", x"eb", x"0a", x"bd",
    x"07", x"04", x"fd", x"fb", x"f8", x"fb", x"01", x"00",
    x"04", x"ff", x"ff", x"fb", x"ff", x"fd", x"fc", x"fb",
    x"00", x"ff", x"36", x"24", x"64", x"35", x"f6", x"37",
    x"78", x"42", x"35", x"29", x"29", x"15", x"24", x"2a",
    x"ce", x"fa", x"1f", x"b5", x"de", x"9f", x"d9", x"c8",
    x"da", x"0a", x"df", x"f3", x"e3", x"07", x"c4", x"04",
    x"13", x"e1", x"db", x"fe", x"de", x"0a", x"c7", x"f1",
    x"d5", x"ac", x"ee", x"f3", x"a1", x"c6", x"f8", x"e0",
    x"1e", x"31", x"32", x"17", x"0b", x"21", x"9e", x"c0",
    x"13", x"27", x"f0", x"13", x"2d", x"fd", x"e0", x"f7",
    x"f8", x"9b", x"17", x"f9", x"d9", x"f4", x"35", x"e4",
    x"0b", x"5f", x"36", x"01", x"e2", x"f3", x"26", x"01",
    x"f3", x"f7", x"f9", x"ec", x"02", x"0f", x"fa", x"04",
    x"df", x"a3", x"ef", x"b4", x"20", x"2d", x"48", x"20",
    x"05", x"26", x"c8", x"16", x"39", x"2d", x"26", x"23",
    x"0b", x"09", x"1b", x"c2", x"fb", x"29", x"01", x"2e",
    x"0f", x"12", x"06", x"f0", x"0d", x"3d", x"ea", x"05",
    x"2b", x"28", x"16", x"fc", x"dd", x"26", x"15", x"fd",
    x"f1", x"0b", x"26", x"04", x"38", x"3b", x"32", x"50",
    x"65", x"10", x"13", x"dd", x"f2", x"24", x"22", x"e2",
    x"01", x"26", x"e5", x"ba", x"ae", x"36", x"39", x"20",
    x"fd", x"fb", x"31", x"f5", x"dd", x"fe", x"35", x"31",
    x"0b", x"ad", x"82", x"c4", x"14", x"14", x"b7", x"43",
    x"f9", x"08", x"e7", x"01", x"f7", x"06", x"f2", x"af",
    x"d9", x"0a", x"ea", x"ec", x"40", x"58", x"ce", x"1a",
    x"17", x"16", x"30", x"57", x"1c", x"03", x"e1", x"07",
    x"44", x"05", x"c8", x"11", x"4a", x"fc", x"13", x"44",
    x"c3", x"eb", x"e8", x"98", x"a8", x"e4", x"11", x"09",
    x"4d", x"f6", x"0a", x"e8", x"38", x"ff", x"c6", x"b8",
    x"bc", x"02", x"2c", x"4b", x"1a", x"41", x"06", x"0e",
    x"15", x"1e", x"00", x"f6", x"fd", x"29", x"c8", x"3d",
    x"08", x"ee", x"3f", x"2a", x"10", x"d8", x"79", x"e8",
    x"fb", x"e7", x"06", x"13", x"06", x"f8", x"fd", x"0e",
    x"04", x"23", x"50", x"f1", x"f9", x"0d", x"f1", x"1d",
    x"22", x"bb", x"c1", x"ff", x"fb", x"e2", x"28", x"17",
    x"ca", x"03", x"ff", x"0d", x"0e", x"fb", x"f5", x"fb",
    x"ea", x"0a", x"ef", x"fe", x"f5", x"e5", x"25", x"fd",
    x"c3", x"05", x"02", x"02", x"fd", x"03", x"02", x"fc",
    x"02", x"04", x"e8", x"f2", x"e7", x"bb", x"ac", x"92",
    x"26", x"18", x"4a", x"03", x"17", x"f7", x"0e", x"18",
    x"f1", x"02", x"42", x"27", x"25", x"49", x"4d", x"12",
    x"27", x"12", x"cf", x"bb", x"a9", x"00", x"fb", x"ca",
    x"15", x"df", x"dc", x"3b", x"41", x"21", x"05", x"3a",
    x"15", x"17", x"0c", x"03", x"27", x"15", x"2a", x"f4",
    x"dd", x"b3", x"e0", x"d1", x"af", x"07", x"ec", x"07",
    x"1f", x"05", x"2c", x"45", x"1c", x"13", x"23", x"17",
    x"05", x"30", x"15", x"0d", x"04", x"1d", x"0a", x"09",
    x"ea", x"b8", x"dd", x"11", x"f2", x"e6", x"ec", x"01",
    x"5f", x"42", x"43", x"02", x"03", x"07", x"fa", x"f3",
    x"06", x"f8", x"00", x"fe", x"09", x"f7", x"0b", x"ec",
    x"c5", x"cc", x"1f", x"dd", x"d9", x"18", x"ef", x"ee",
    x"0c", x"f9", x"2c", x"01", x"ba", x"95", x"c6", x"ed",
    x"ed", x"03", x"de", x"f3", x"c3", x"e1", x"f6", x"e4",
    x"c2", x"aa", x"c3", x"de", x"ec", x"fd", x"04", x"f1",
    x"12", x"01", x"1d", x"c1", x"da", x"0b", x"2b", x"1b",
    x"ed", x"e3", x"f6", x"e5", x"00", x"df", x"ba", x"b4",
    x"b4", x"ce", x"d7", x"f7", x"ee", x"0d", x"5e", x"26",
    x"e0", x"28", x"13", x"0f", x"e4", x"23", x"df", x"16",
    x"fc", x"ee", x"df", x"ea", x"05", x"fb", x"f9", x"04",
    x"f7", x"fa", x"00", x"01", x"0f", x"73", x"1e", x"05",
    x"30", x"24", x"ea", x"e5", x"be", x"c4", x"66", x"f0",
    x"0a", x"1b", x"f8", x"f8", x"29", x"d2", x"e2", x"e5",
    x"1b", x"45", x"e0", x"eb", x"0e", x"0f", x"09", x"fe",
    x"00", x"ff", x"fd", x"03", x"fd", x"01", x"fc", x"fb",
    x"01", x"ca", x"da", x"f7", x"d5", x"e8", x"d4", x"d0",
    x"16", x"c7", x"02", x"10", x"1c", x"f6", x"fe", x"e6",
    x"20", x"10", x"16", x"10", x"db", x"10", x"f6", x"ee",
    x"1d", x"2d", x"d9", x"c6", x"07", x"67", x"55", x"2e",
    x"29", x"24", x"3d", x"2d", x"ea", x"a0", x"9e", x"22",
    x"ea", x"0b", x"15", x"12", x"f5", x"05", x"3d", x"36",
    x"0d", x"f3", x"ce", x"0c", x"f8", x"ec", x"03", x"fc",
    x"00", x"11", x"f8", x"ec", x"aa", x"34", x"5f", x"76",
    x"00", x"ff", x"00", x"06", x"fc", x"07", x"01", x"00",
    x"01", x"03", x"08", x"02", x"05", x"fc", x"fc", x"01",
    x"fd", x"00", x"14", x"c6", x"7f", x"e5", x"d1", x"c1",
    x"05", x"f1", x"fe", x"f1", x"19", x"4b", x"14", x"18",
    x"1b", x"15", x"17", x"e3", x"12", x"2c", x"23", x"0e",
    x"18", x"c6", x"02", x"1b", x"49", x"e0", x"d2", x"c3",
    x"04", x"ee", x"0a", x"31", x"41", x"35", x"0a", x"2f",
    x"39", x"de", x"29", x"fa", x"f2", x"00", x"f0", x"18",
    x"f1", x"13", x"03", x"30", x"28", x"f4", x"21", x"df",
    x"13", x"2e", x"2c", x"19", x"12", x"0d", x"18", x"ec",
    x"b2", x"05", x"fb", x"17", x"d1", x"bd", x"e1", x"f3",
    x"e8", x"d9", x"f3", x"22", x"34", x"0f", x"03", x"02",
    x"2e", x"d5", x"fd", x"d7", x"f2", x"e6", x"68", x"08",
    x"06", x"21", x"22", x"21", x"15", x"f7", x"bf", x"10",
    x"db", x"ad", x"eb", x"e8", x"de", x"0b", x"fc", x"0a",
    x"eb", x"df", x"cb", x"2a", x"c3", x"ca", x"ef", x"d2",
    x"94", x"b6", x"de", x"d7", x"fc", x"26", x"31", x"a3",
    x"b9", x"df", x"29", x"29", x"14", x"fc", x"ee", x"e7",
    x"cc", x"fa", x"15", x"d8", x"ed", x"ec", x"fb", x"e9",
    x"57", x"e1", x"f4", x"29", x"fa", x"ec", x"d4", x"16",
    x"0a", x"08", x"32", x"29", x"3e", x"5b", x"2b", x"1a",
    x"f6", x"0b", x"14", x"01", x"f3", x"08", x"1f", x"01",
    x"10", x"f1", x"07", x"bc", x"07", x"f6", x"56", x"28",
    x"18", x"04", x"12", x"00", x"0a", x"28", x"2d", x"c1",
    x"12", x"f3", x"f6", x"de", x"fb", x"10", x"f1", x"9f",
    x"d4", x"cf", x"c3", x"09", x"db", x"e7", x"32", x"eb",
    x"99", x"0c", x"c3", x"ce", x"e4", x"de", x"01", x"03",
    x"e3", x"cc", x"cd", x"f7", x"09", x"0a", x"17", x"05",
    x"fb", x"39", x"0c", x"f9", x"eb", x"f0", x"ff", x"10",
    x"0d", x"ec", x"2a", x"17", x"2e", x"78", x"42", x"23",
    x"5a", x"50", x"31", x"b7", x"9c", x"f3", x"00", x"b3",
    x"06", x"1f", x"e8", x"0d", x"6b", x"63", x"27", x"ba",
    x"eb", x"e7", x"1b", x"11", x"fc", x"d5", x"4a", x"44",
    x"0b", x"2a", x"50", x"0a", x"00", x"f4", x"43", x"28",
    x"d2", x"e1", x"c9", x"f1", x"ef", x"04", x"11", x"b1",
    x"ed", x"ae", x"b3", x"24", x"23", x"ef", x"17", x"fe",
    x"b5", x"c0", x"8b", x"e6", x"e9", x"be", x"d1", x"d8",
    x"e0", x"ff", x"fc", x"fc", x"00", x"00", x"04", x"04",
    x"01", x"fc", x"3c", x"1a", x"26", x"0c", x"e1", x"8e",
    x"02", x"0f", x"0f", x"f7", x"00", x"5a", x"07", x"23",
    x"10", x"fc", x"e3", x"f3", x"bb", x"ff", x"26", x"c9",
    x"b1", x"34", x"f1", x"e6", x"12", x"36", x"1a", x"20",
    x"13", x"02", x"34", x"e3", x"eb", x"03", x"ca", x"fd",
    x"b8", x"d0", x"e6", x"05", x"f0", x"10", x"0c", x"c7",
    x"e0", x"e8", x"1e", x"2d", x"22", x"24", x"05", x"03",
    x"e7", x"b6", x"c6", x"16", x"f6", x"e8", x"26", x"05",
    x"02", x"14", x"0e", x"11", x"06", x"24", x"3f", x"18",
    x"10", x"16", x"50", x"1b", x"16", x"53", x"17", x"1e",
    x"16", x"e3", x"f7", x"0e", x"07", x"fa", x"0a", x"02",
    x"0a", x"06", x"0c", x"01", x"0b", x"e2", x"f1", x"d6",
    x"f1", x"da", x"b6", x"f2", x"dd", x"e0", x"09", x"bf",
    x"17", x"16", x"e4", x"3d", x"1f", x"0c", x"61", x"13",
    x"18", x"3a", x"0b", x"0b", x"07", x"02", x"06", x"b0",
    x"97", x"03", x"c2", x"ef", x"0e", x"1a", x"19", x"10",
    x"95", x"8b", x"e9", x"09", x"25", x"47", x"0e", x"01",
    x"da", x"1f", x"13", x"19", x"2e", x"03", x"0d", x"17",
    x"f8", x"16", x"eb", x"e8", x"24", x"a3", x"c6", x"c3",
    x"e7", x"d1", x"c7", x"c5", x"09", x"1b", x"03", x"01",
    x"fd", x"3d", x"f5", x"fc", x"05", x"ff", x"0c", x"03",
    x"fd", x"02", x"01", x"03", x"06", x"6d", x"6d", x"58",
    x"0b", x"09", x"2f", x"ea", x"f2", x"18", x"49", x"1c",
    x"ff", x"46", x"43", x"f2", x"21", x"00", x"06", x"d6",
    x"ad", x"e6", x"d6", x"3d", x"02", x"36", x"12", x"0a",
    x"fb", x"fe", x"03", x"fe", x"01", x"fd", x"ff", x"01",
    x"fc", x"f1", x"ef", x"11", x"37", x"2d", x"1c", x"f8",
    x"16", x"09", x"c7", x"82", x"0a", x"9d", x"d7", x"11",
    x"e1", x"16", x"e8", x"76", x"4e", x"27", x"55", x"26",
    x"10", x"13", x"ed", x"e5", x"4c", x"13", x"18", x"1e",
    x"dd", x"13", x"eb", x"c3", x"f8", x"bc", x"c1", x"b2",
    x"be", x"0d", x"37", x"cf", x"00", x"40", x"5c", x"31",
    x"b6", x"69", x"14", x"b2", x"05", x"f8", x"0b", x"74",
    x"39", x"19", x"50", x"16", x"17", x"f8", x"06", x"19",
    x"fd", x"02", x"0b", x"04", x"04", x"01", x"ff", x"04",
    x"fa", x"02", x"05", x"02", x"fe", x"02", x"03", x"07",
    x"07", x"07", x"3c", x"dc", x"cb", x"d9", x"da", x"bd",
    x"0a", x"fe", x"f3", x"47", x"ed", x"1d", x"2a", x"28",
    x"16", x"15", x"fd", x"e6", x"5e", x"75", x"28", x"4c",
    x"39", x"24", x"ea", x"e6", x"20", x"bb", x"dc", x"04",
    x"16", x"f6", x"d3", x"1d", x"04", x"b6", x"ec", x"b2",
    x"d4", x"31", x"de", x"e0", x"e8", x"e4", x"e6", x"c3",
    x"59", x"87", x"ec", x"b3", x"cf", x"3d", x"0c", x"0a",
    x"d4", x"d8", x"bb", x"17", x"d4", x"fe", x"3f", x"f6",
    x"fd", x"d2", x"f0", x"50", x"4e", x"2d", x"01", x"57",
    x"0f", x"1d", x"26", x"13", x"ef", x"b3", x"fa", x"0f",
    x"fa", x"12", x"17", x"58", x"1b", x"06", x"14", x"ea",
    x"f8", x"f6", x"e7", x"19", x"d5", x"e9", x"e7", x"b1",
    x"f0", x"fa", x"33", x"1e", x"1e", x"ce", x"fd", x"f5",
    x"09", x"19", x"00", x"05", x"08", x"ef", x"bd", x"b5",
    x"c9", x"15", x"f5", x"da", x"fd", x"0b", x"ef", x"6e",
    x"25", x"ae", x"c6", x"06", x"b6", x"e1", x"12", x"ed",
    x"fd", x"fd", x"04", x"04", x"00", x"fb", x"00", x"fc",
    x"01", x"ff", x"fd", x"01", x"ff", x"fa", x"fb", x"fd",
    x"fd", x"fc", x"ff", x"04", x"00", x"fd", x"04", x"fe",
    x"04", x"ff", x"fb", x"fe", x"f8", x"fc", x"ff", x"fc",
    x"fe", x"fc", x"fb", x"f8", x"fc", x"ff", x"fe", x"02",
    x"fb", x"04", x"01", x"01", x"01", x"fa", x"02", x"fe",
    x"ff", x"fc", x"04", x"fe", x"fa", x"04", x"03", x"fe",
    x"00", x"ff", x"fd", x"00", x"fe", x"fa", x"02", x"fb",
    x"fe", x"fc", x"00", x"01", x"fb", x"ff", x"00", x"02",
    x"04", x"03", x"01", x"02", x"fd", x"03", x"00", x"fb",
    x"fd", x"fc", x"fd", x"ff", x"00", x"fb", x"fc", x"f9",
    x"00", x"f9", x"03", x"fc", x"02", x"fc", x"fc", x"fe",
    x"02", x"02", x"01", x"fe", x"fd", x"02", x"03", x"fb",
    x"fc", x"03", x"fc", x"03", x"fc", x"fd", x"02", x"fe",
    x"04", x"fc", x"02", x"01", x"fb", x"fd", x"fd", x"06",
    x"f6", x"fd", x"fc", x"fd", x"fd", x"fd", x"04", x"fa",
    x"04", x"02", x"00", x"fa", x"fd", x"fd", x"fb", x"fc",
    x"ff", x"fa", x"f8", x"fe", x"00", x"03", x"fd", x"fd",
    x"00", x"01", x"fa", x"fa", x"fa", x"01", x"ff", x"01",
    x"ff", x"00", x"ff", x"03", x"00", x"fe", x"02", x"fd",
    x"fb", x"00", x"05", x"01", x"fc", x"00", x"fb", x"04",
    x"fb", x"fb", x"02", x"01", x"01", x"00", x"fa", x"fd",
    x"04", x"ff", x"fb", x"fa", x"fe", x"00", x"00", x"02",
    x"03", x"04", x"f9", x"ff", x"02", x"04", x"00", x"fa",
    x"00", x"fd", x"ff", x"03", x"f9", x"00", x"fe", x"fe",
    x"03", x"ff", x"03", x"00", x"fc", x"ff", x"04", x"fd",
    x"01", x"fd", x"ff", x"fc", x"01", x"ff", x"00", x"fe",
    x"02", x"fc", x"fb", x"fe", x"fd", x"01", x"04", x"f8",
    x"f8", x"ff", x"03", x"ff", x"fa", x"fe", x"ff", x"fd",
    x"01", x"fb", x"00", x"fd", x"fb", x"fd", x"ff", x"fc",
    x"fd", x"f9", x"fd", x"fe", x"04", x"00", x"04", x"02",
    x"ff", x"00", x"fe", x"05", x"fd", x"01", x"fc", x"fa",
    x"fa", x"fb", x"fb", x"02", x"fd", x"03", x"02", x"00",
    x"f8", x"02", x"00", x"f9", x"03", x"01", x"fd", x"ff",
    x"fd", x"fa", x"fa", x"f7", x"fe", x"00", x"fe", x"03",
    x"02", x"02", x"03", x"fb", x"ff", x"fe", x"fb", x"03",
    x"fc", x"fa", x"01", x"fd", x"f9", x"fc", x"f9", x"ff",
    x"fd", x"fc", x"01", x"00", x"04", x"fc", x"fa", x"fd",
    x"f7", x"00", x"ff", x"fb", x"00", x"fd", x"04", x"fe",
    x"02", x"ff", x"01", x"03", x"fd", x"fd", x"00", x"f6",
    x"00", x"fe", x"f8", x"03", x"02", x"04", x"fe", x"02",
    x"03", x"fe", x"04", x"00", x"ff", x"ff", x"ff", x"03",
    x"04", x"03", x"fb", x"03", x"f6", x"03", x"fb", x"fe",
    x"03", x"02", x"fc", x"04", x"fb", x"fc", x"fa", x"00",
    x"fb", x"01", x"fd", x"04", x"fb", x"f6", x"fc", x"fb",
    x"fb", x"04", x"04", x"fe", x"04", x"fe", x"ff", x"fe",
    x"fb", x"03", x"03", x"04", x"fc", x"00", x"fd", x"01",
    x"04", x"00", x"fa", x"fc", x"02", x"fc", x"02", x"fe",
    x"fb", x"ff", x"ff", x"02", x"fb", x"04", x"fb", x"fc",
    x"04", x"fd", x"fd", x"fd", x"fa", x"fb", x"00", x"01",
    x"fd", x"fb", x"00", x"f9", x"fe", x"fe", x"ff", x"02",
    x"fa", x"fc", x"01", x"fe", x"01", x"fe", x"fe", x"00",
    x"02", x"fa", x"fa", x"fa", x"fb", x"fc", x"fb", x"ff",
    x"fb", x"fd", x"fe", x"01", x"01", x"fa", x"fb", x"fc",
    x"ff", x"ff", x"04", x"04", x"fd", x"fe", x"00", x"00",
    x"00", x"fb", x"03", x"00", x"03", x"05", x"fe", x"00",
    x"03", x"fd", x"02", x"fb", x"fc", x"fc", x"fd", x"ff",
    x"fd", x"f8", x"ff", x"02", x"fd", x"01", x"fe", x"03",
    x"fd", x"f8", x"fb", x"04", x"04", x"fb", x"02", x"ff",
    x"fb", x"fe", x"fb", x"f6", x"04", x"02", x"02", x"fd",
    x"fb", x"f9", x"fb", x"fb", x"02", x"fe", x"fb", x"01",
    x"02", x"fc", x"01", x"fd", x"fc", x"fd", x"fb", x"02",
    x"03", x"ff", x"01", x"f7", x"fa", x"fa", x"fe", x"01",
    x"fd", x"00", x"fb", x"01", x"fd", x"fe", x"02", x"03",
    x"fe", x"fc", x"ff", x"04", x"02", x"f7", x"04", x"fd",
    x"fe", x"00", x"01", x"01", x"fc", x"00", x"fb", x"fc",
    x"fc", x"fd", x"fb", x"02", x"01", x"00", x"00", x"f7",
    x"f9", x"fe", x"00", x"fd", x"fe", x"03", x"02", x"00",
    x"fc", x"00", x"02", x"fc", x"fd", x"fb", x"01", x"fc",
    x"fd", x"fa", x"ff", x"f7", x"fd", x"fe", x"05", x"fd",
    x"fe", x"00", x"00", x"fb", x"02", x"01", x"fe", x"03",
    x"ff", x"ff", x"fd", x"01", x"fb", x"fd", x"ff", x"00",
    x"fb", x"fe", x"02", x"fc", x"fb", x"fe", x"fc", x"f7",
    x"08", x"03", x"02", x"f6", x"03", x"fa", x"00", x"ff",
    x"fb", x"fd", x"ff", x"fb", x"ff", x"04", x"fe", x"fb",
    x"fd", x"f8", x"ff", x"fd", x"fc", x"fa", x"f8", x"01",
    x"fb", x"fc", x"03", x"fc", x"04", x"00", x"fb", x"04",
    x"03", x"fb", x"fe", x"fd", x"fe", x"fc", x"fd", x"f9",
    x"fb", x"03", x"f7", x"fd", x"f7", x"00", x"04", x"ff",
    x"fb", x"03", x"fa", x"f9", x"04", x"f9", x"f5", x"02",
    x"fc", x"02", x"fd", x"fa", x"fe", x"00", x"fb", x"ff",
    x"03", x"fb", x"01", x"ff", x"fd", x"03", x"fe", x"fd",
    x"fd", x"fb", x"f6", x"f4", x"fc", x"f8", x"03", x"fc",
    x"f6", x"fc", x"fe", x"00", x"f7", x"fc", x"04", x"02",
    x"fe", x"00", x"fc", x"ff", x"04", x"fb", x"04", x"01",
    x"f7", x"01", x"04", x"f7", x"01", x"ff", x"fd", x"00",
    x"04", x"fa", x"04", x"fb", x"f6", x"fe", x"fd", x"03",
    x"04", x"ff", x"02", x"fd", x"01", x"f9", x"02", x"f9",
    x"01", x"fe", x"fe", x"fd", x"fa", x"fe", x"fb", x"00",
    x"fc", x"f9", x"f7", x"fc", x"fb", x"f7", x"fb", x"02",
    x"02", x"fb", x"fd", x"fb", x"01", x"f8", x"03", x"00",
    x"fa", x"fe", x"04", x"00", x"03", x"01", x"ff", x"04",
    x"04", x"01", x"fe", x"fd", x"fc", x"fc", x"01", x"f6",
    x"00", x"fc", x"fb", x"fa", x"fd", x"fc", x"01", x"06",
    x"fa", x"fd", x"fb", x"f9", x"f9", x"00", x"f7", x"fc",
    x"fe", x"02", x"fa", x"fd", x"00", x"01", x"fa", x"00",
    x"03", x"04", x"f6", x"00", x"fb", x"fb", x"fe", x"03",
    x"f9", x"01", x"fd", x"01", x"f9", x"f6", x"ff", x"04",
    x"00", x"f7", x"fa", x"fd", x"ff", x"00", x"ff", x"f7",
    x"fd", x"01", x"fb", x"00", x"03", x"fd", x"04", x"01",
    x"fe", x"01", x"ff", x"fd", x"04", x"00", x"fe", x"fe",
    x"00", x"f7", x"fd", x"f8", x"fa", x"03", x"01", x"fe",
    x"fb", x"01", x"fb", x"01", x"00", x"00", x"04", x"fc",
    x"03", x"01", x"fd", x"fc", x"fa", x"fb", x"fc", x"fd",
    x"fb", x"00", x"fd", x"f7", x"f5", x"ff", x"fb", x"ff",
    x"f8", x"fe", x"fe", x"02", x"fa", x"f9", x"04", x"fc",
    x"fd", x"fe", x"02", x"03", x"00", x"fe", x"03", x"fc",
    x"00", x"fa", x"fb", x"fd", x"fc", x"fb", x"fa", x"fc",
    x"fa", x"f9", x"fc", x"ff", x"fa", x"fd", x"00", x"fc",
    x"00", x"f7", x"fe", x"f7", x"00", x"f8", x"02", x"f9",
    x"f7", x"fd", x"fb", x"00", x"f8", x"fa", x"ff", x"fe",
    x"fd", x"f8", x"04", x"00", x"f9", x"fd", x"fd", x"fd",
    x"fa", x"fa", x"fa", x"fb", x"ff", x"00", x"05", x"01",
    x"fd", x"fe", x"ff", x"02", x"01", x"02", x"fe", x"fe",
    x"fa", x"ff", x"00", x"01", x"fc", x"06", x"fe", x"02",
    x"fe", x"04", x"fc", x"01", x"04", x"ff", x"fb", x"f8",
    x"fb", x"ff", x"fd", x"fe", x"f9", x"ff", x"00", x"fa",
    x"fe", x"00", x"00", x"03", x"fb", x"05", x"03", x"ff",
    x"01", x"00", x"fd", x"fa", x"fb", x"fd", x"fa", x"04",
    x"fd", x"00", x"fc", x"00", x"f8", x"fd", x"f8", x"ff",
    x"fe", x"fb", x"fc", x"fa", x"ff", x"fb", x"fb", x"fe",
    x"f9", x"00", x"fd", x"fc", x"00", x"00", x"02", x"02",
    x"ff", x"03", x"01", x"fe", x"01", x"fb", x"04", x"fd",
    x"fb", x"ff", x"fa", x"01", x"f9", x"f8", x"fb", x"fb",
    x"fe", x"fb", x"00", x"f9", x"02", x"fb", x"01", x"ff",
    x"f7", x"fc", x"ff", x"04", x"fd", x"fb", x"fb", x"f9",
    x"02", x"fe", x"02", x"01", x"fe", x"01", x"ff", x"fe",
    x"ff", x"ff", x"05", x"00", x"04", x"01", x"fb", x"02",
    x"fd", x"01", x"fd", x"fa", x"fd", x"fc", x"ff", x"02",
    x"f9", x"fc", x"06", x"ff", x"fe", x"fb", x"fe", x"fe",
    x"fd", x"fa", x"fc", x"fe", x"fb", x"fd", x"f7", x"fc",
    x"fa", x"fa", x"fa", x"03", x"fe", x"03", x"fc", x"fc",
    x"f9", x"f9", x"f7", x"fd", x"fc", x"f9", x"fd", x"01",
    x"03", x"00", x"fd", x"fc", x"fb", x"ff", x"fe", x"fa",
    x"01", x"00", x"fc", x"ff", x"fa", x"00", x"fd", x"f8",
    x"fe", x"ff", x"ff", x"fc", x"00", x"00", x"f8", x"04",
    x"fb", x"fa", x"fa", x"f8", x"fa", x"fa", x"f6", x"fc",
    x"ff", x"fa", x"00", x"00", x"f8", x"fb", x"fb", x"fd",
    x"02", x"fb", x"01", x"03", x"01", x"f9", x"fe", x"fe",
    x"ff", x"fb", x"f9", x"f7", x"ff", x"fb", x"fa", x"fa",
    x"04", x"01", x"03", x"01", x"fb", x"fa", x"ff", x"fb",
    x"01", x"fb", x"ff", x"fb", x"03", x"fb", x"fe", x"fd",
    x"fc", x"00", x"fc", x"fa", x"fa", x"fe", x"f5", x"02",
    x"fa", x"f8", x"03", x"fb", x"f9", x"ff", x"f8", x"00",
    x"01", x"fd", x"fa", x"fe", x"fc", x"02", x"fa", x"ff",
    x"fb", x"01", x"ff", x"fe", x"fb", x"fe", x"f7", x"04",
    x"fa", x"fb", x"01", x"fb", x"02", x"00", x"ff", x"ff",
    x"00", x"fe", x"00", x"f4", x"fe", x"02", x"fa", x"fb",
    x"00", x"fe", x"f5", x"02", x"fd", x"fa", x"fc", x"04",
    x"fb", x"ff", x"ff", x"fd", x"03", x"fe", x"02", x"fe",
    x"00", x"fb", x"f9", x"fe", x"04", x"fb", x"fc", x"00",
    x"fc", x"00", x"fd", x"03", x"01", x"fc", x"fe", x"fb",
    x"04", x"ff", x"ff", x"f9", x"04", x"fe", x"fe", x"fc",
    x"ff", x"fe", x"02", x"fe", x"fa", x"fc", x"01", x"fa",
    x"fd", x"fc", x"fe", x"fe", x"fb", x"01", x"00", x"fd",
    x"ff", x"04", x"fb", x"04", x"fc", x"fa", x"03", x"f9",
    x"fd", x"fe", x"fc", x"fa", x"03", x"ff", x"fa", x"fd",
    x"fb", x"fb", x"01", x"f8", x"fb", x"f8", x"fb", x"03",
    x"f8", x"fb", x"fd", x"01", x"01", x"f9", x"fa", x"fc",
    x"fa", x"fd", x"03", x"fa", x"fb", x"ff", x"ff", x"fd",
    x"fc", x"fe", x"fc", x"fb", x"02", x"fd", x"ff", x"fe",
    x"03", x"fc", x"fa", x"04", x"fd", x"00", x"fa", x"01",
    x"fa", x"fb", x"03", x"fe", x"f7", x"fd", x"fb", x"fa",
    x"fc", x"03", x"01", x"fc", x"fc", x"00", x"00", x"fd",
    x"00", x"02", x"03", x"03", x"00", x"fa", x"fb", x"ff",
    x"00", x"fa", x"00", x"fe", x"fc", x"fe", x"01", x"f9",
    x"fa", x"fc", x"03", x"fa", x"02", x"fa", x"00", x"fd",
    x"fd", x"fa", x"ff", x"fb", x"fd", x"04", x"01", x"f5",
    x"04", x"00", x"f9", x"fd", x"ff", x"03", x"02", x"ff",
    x"fe", x"fb", x"f7", x"00", x"fe", x"fb", x"01", x"f9",
    x"fd", x"fe", x"fe", x"fc", x"fb", x"fd", x"02", x"fd",
    x"02", x"ff", x"01", x"fe", x"fd", x"01", x"03", x"fb",
    x"f8", x"fc", x"00", x"fd", x"01", x"fe", x"fb", x"fb",
    x"ff", x"00", x"fc", x"fa", x"f8", x"01", x"fe", x"ff",
    x"fc", x"00", x"04", x"fb", x"fb", x"04", x"ff", x"01",
    x"02", x"ff", x"01", x"fd", x"fa", x"fa", x"02", x"00",
    x"fe", x"ff", x"fd", x"00", x"ff", x"02", x"fc", x"02",
    x"fc", x"ff", x"fd", x"01", x"01", x"02", x"ff", x"03",
    x"ff", x"03", x"fd", x"fd", x"02", x"04", x"00", x"fe",
    x"fd", x"f9", x"ff", x"ff", x"fe", x"01", x"fe", x"01",
    x"02", x"f8", x"f9", x"fd", x"00", x"ff", x"f9", x"02",
    x"ff", x"ff", x"fe", x"02", x"fb", x"f9", x"00", x"fd",
    x"f5", x"01", x"00", x"00", x"ff", x"01", x"ff", x"fb",
    x"01", x"03", x"fb", x"02", x"fb", x"04", x"00", x"fa",
    x"fc", x"03", x"fd", x"f9", x"fd", x"fd", x"05", x"fe",
    x"ff", x"04", x"05", x"01", x"01", x"fa", x"00", x"fe",
    x"04", x"ff", x"fa", x"03", x"fe", x"03", x"00", x"fe",
    x"fa", x"fc", x"fb", x"f9", x"fc", x"fc", x"f6", x"ff",
    x"ff", x"f7", x"fe", x"01", x"fc", x"02", x"f9", x"f9",
    x"01", x"fe", x"fd", x"fd", x"06", x"fd", x"fd", x"05",
    x"ff", x"ff", x"fc", x"01", x"00", x"ff", x"f7", x"02",
    x"00", x"fe", x"00", x"fe", x"fe", x"ff", x"fc", x"fd",
    x"ff", x"02", x"02", x"fb", x"02", x"f7", x"fc", x"fb",
    x"01", x"fe", x"fe", x"fd", x"05", x"02", x"03", x"02",
    x"03", x"fe", x"00", x"ff", x"fd", x"f8", x"fd", x"fb",
    x"fb", x"02", x"01", x"fe", x"fa", x"fb", x"fe", x"fb",
    x"f8", x"00", x"01", x"ff", x"03", x"fb", x"fe", x"fb",
    x"fd", x"fa", x"fb", x"f9", x"04", x"02", x"01", x"01",
    x"00", x"fe", x"fc", x"fc", x"01", x"fc", x"fe", x"05",
    x"ff", x"02", x"ff", x"fb", x"fb", x"02", x"fe", x"02",
    x"fc", x"02", x"02", x"fd", x"00", x"ff", x"f9", x"03",
    x"05", x"fe", x"ff", x"01", x"03", x"fb", x"00", x"01",
    x"03", x"00", x"01", x"02", x"ff", x"fe", x"fc", x"03",
    x"fa", x"fa", x"00", x"03", x"00", x"00", x"fa", x"f5",
    x"00", x"fc", x"fb", x"04", x"fb", x"fb", x"01", x"f8",
    x"fb", x"f9", x"f8", x"fc", x"03", x"fb", x"fe", x"02",
    x"01", x"fb", x"02", x"fb", x"ff", x"04", x"02", x"00",
    x"fb", x"fd", x"04", x"ff", x"02", x"fa", x"00", x"00",
    x"ff", x"fc", x"fb", x"f8", x"01", x"fc", x"fe", x"04",
    x"03", x"01", x"00", x"fd", x"fc", x"fa", x"03", x"fd",
    x"fc", x"ff", x"ff", x"f8", x"fb", x"00", x"fe", x"fe",
    x"fd", x"00", x"fe", x"04", x"fb", x"00", x"fd", x"04",
    x"fd", x"f8", x"fc", x"02", x"fd", x"04", x"fc", x"01",
    x"fa", x"ff", x"f8", x"fe", x"fe", x"fd", x"02", x"fa",
    x"f9", x"fc", x"f8", x"03", x"fe", x"fd", x"ff", x"fe",
    x"02", x"01", x"fd", x"fd", x"fe", x"03", x"01", x"fa",
    x"dd", x"d8", x"24", x"f1", x"e6", x"f6", x"f8", x"f3",
    x"d3", x"dd", x"c9", x"0c", x"d8", x"e7", x"04", x"ee",
    x"1d", x"18", x"d5", x"0a", x"e3", x"04", x"fb", x"0b",
    x"4c", x"14", x"17", x"32", x"2f", x"00", x"f2", x"b8",
    x"b8", x"e1", x"fd", x"df", x"d2", x"c7", x"ca", x"e2",
    x"b6", x"d9", x"2e", x"33", x"5b", x"3f", x"17", x"f4",
    x"10", x"fc", x"3a", x"d3", x"07", x"2c", x"26", x"dd",
    x"1b", x"f9", x"e7", x"ef", x"e3", x"a5", x"a5", x"d0",
    x"a6", x"f2", x"29", x"28", x"10", x"e4", x"d3", x"c2",
    x"c9", x"e4", x"fe", x"30", x"1f", x"38", x"04", x"e3",
    x"0a", x"0f", x"35", x"4e", x"49", x"0a", x"22", x"f4",
    x"e7", x"df", x"de", x"a9", x"cf", x"f9", x"ab", x"ab",
    x"45", x"ca", x"db", x"f3", x"f4", x"16", x"20", x"30",
    x"18", x"22", x"d0", x"c8", x"26", x"f2", x"fe", x"ef",
    x"3e", x"26", x"dd", x"ff", x"fe", x"a5", x"85", x"a1",
    x"e3", x"f7", x"a2", x"33", x"f9", x"40", x"a9", x"d8",
    x"f4", x"0a", x"01", x"17", x"28", x"2a", x"0a", x"ff",
    x"19", x"3a", x"29", x"2c", x"4c", x"4e", x"25", x"ee",
    x"2e", x"df", x"d3", x"08", x"f9", x"12", x"f9", x"fb",
    x"ea", x"01", x"ff", x"ff", x"fc", x"01", x"00", x"04",
    x"03", x"03", x"e1", x"81", x"ab", x"ff", x"a2", x"0c",
    x"f4", x"ce", x"e0", x"e6", x"03", x"e9", x"fe", x"ec",
    x"e2", x"04", x"23", x"f5", x"ac", x"a5", x"ab", x"31",
    x"02", x"f2", x"fc", x"e1", x"cf", x"d3", x"1d", x"2a",
    x"ec", x"0a", x"ff", x"e9", x"04", x"f8", x"df", x"f0",
    x"f9", x"f6", x"d2", x"e2", x"0b", x"f6", x"c0", x"bf",
    x"ef", x"fd", x"cd", x"fb", x"0c", x"30", x"25", x"12",
    x"ce", x"99", x"d7", x"33", x"a0", x"b7", x"eb", x"5d",
    x"2d", x"e5", x"c9", x"fc", x"3d", x"30", x"fc", x"48",
    x"53", x"2c", x"1e", x"f7", x"0d", x"2d", x"10", x"1d",
    x"15", x"1c", x"23", x"00", x"02", x"00", x"fa", x"ff",
    x"06", x"06", x"fa", x"fe", x"d9", x"0b", x"03", x"ee",
    x"06", x"fb", x"17", x"1c", x"d3", x"1b", x"30", x"ec",
    x"f6", x"f8", x"06", x"e0", x"c4", x"fa", x"1d", x"d8",
    x"f8", x"0a", x"ef", x"e3", x"1a", x"fc", x"ff", x"f5",
    x"ed", x"fc", x"21", x"25", x"31", x"f8", x"ff", x"fe",
    x"b8", x"76", x"db", x"4d", x"65", x"24", x"04", x"fe",
    x"04", x"f7", x"ac", x"f7", x"35", x"28", x"e0", x"09",
    x"cd", x"e9", x"ca", x"04", x"12", x"2d", x"1c", x"41",
    x"2b", x"0c", x"33", x"c2", x"f5", x"f3", x"fb", x"09",
    x"ef", x"a1", x"f1", x"d4", x"0d", x"01", x"03", x"0e",
    x"0c", x"10", x"10", x"11", x"04", x"cd", x"d7", x"c9",
    x"ec", x"ba", x"b5", x"16", x"f2", x"b9", x"07", x"c5",
    x"fe", x"d8", x"e7", x"07", x"6c", x"0c", x"25", x"f0",
    x"e9", x"19", x"1e", x"e5", x"bf", x"0f", x"e9", x"f6",
    x"ff", x"ff", x"fb", x"fb", x"04", x"05", x"ff", x"fb",
    x"fc", x"f9", x"e0", x"bf", x"de", x"e7", x"ed", x"0a",
    x"09", x"e0", x"ac", x"b6", x"b1", x"f9", x"d0", x"ec",
    x"ac", x"93", x"ce", x"32", x"eb", x"fa", x"fc", x"c2",
    x"d2", x"51", x"f3", x"fe", x"3b", x"fc", x"b9", x"10",
    x"c7", x"71", x"0e", x"1b", x"18", x"f7", x"e7", x"d5",
    x"13", x"06", x"1b", x"13", x"1b", x"f5", x"cb", x"c7",
    x"ad", x"c8", x"0d", x"1f", x"2f", x"1a", x"27", x"bf",
    x"54", x"21", x"f8", x"11", x"30", x"46", x"34", x"61",
    x"fc", x"fd", x"fe", x"05", x"fc", x"03", x"fd", x"fc",
    x"ff", x"01", x"01", x"fc", x"fe", x"01", x"01", x"fd",
    x"fc", x"03", x"d2", x"e1", x"e9", x"c5", x"05", x"ec",
    x"3a", x"42", x"32", x"b3", x"9d", x"a4", x"d7", x"c9",
    x"93", x"fb", x"03", x"17", x"ea", x"df", x"f1", x"fa",
    x"17", x"1c", x"ec", x"de", x"0c", x"e8", x"0d", x"fc",
    x"05", x"f7", x"12", x"f4", x"f6", x"bf", x"49", x"e1",
    x"01", x"69", x"3b", x"1f", x"f0", x"d8", x"19", x"ba",
    x"95", x"bb", x"f7", x"ed", x"d2", x"dd", x"e2", x"cd",
    x"ce", x"9a", x"d1", x"ef", x"a6", x"e2", x"d5", x"af",
    x"e4", x"50", x"0b", x"00", x"11", x"16", x"10", x"f5",
    x"f4", x"13", x"cb", x"03", x"e7", x"da", x"0c", x"08",
    x"36", x"22", x"f2", x"1a", x"05", x"ef", x"0c", x"16",
    x"16", x"fe", x"e3", x"10", x"f5", x"34", x"b8", x"0c",
    x"f5", x"e8", x"0f", x"db", x"e2", x"ce", x"05", x"02",
    x"ea", x"1d", x"0b", x"04", x"f1", x"cc", x"de", x"2a",
    x"dc", x"03", x"f0", x"03", x"16", x"ec", x"33", x"c2",
    x"e3", x"14", x"36", x"1f", x"2c", x"d7", x"1f", x"5f",
    x"e8", x"20", x"20", x"c8", x"c9", x"0d", x"a3", x"bd",
    x"2a", x"49", x"07", x"eb", x"c9", x"dc", x"01", x"85",
    x"f3", x"42", x"df", x"22", x"2f", x"15", x"1a", x"2a",
    x"26", x"15", x"46", x"06", x"01", x"1c", x"01", x"f9",
    x"f6", x"bf", x"b6", x"fd", x"03", x"16", x"2b", x"1f",
    x"30", x"23", x"11", x"05", x"de", x"11", x"20", x"1a",
    x"d7", x"07", x"27", x"a7", x"d2", x"f3", x"a9", x"8d",
    x"82", x"d2", x"0c", x"16", x"fd", x"26", x"2a", x"5f",
    x"24", x"0d", x"f8", x"f7", x"c7", x"f2", x"fc", x"df",
    x"17", x"3c", x"52", x"16", x"e7", x"0d", x"f1", x"f6",
    x"1c", x"13", x"1e", x"2e", x"4e", x"3a", x"44", x"5e",
    x"20", x"1b", x"33", x"15", x"11", x"66", x"f3", x"19",
    x"2e", x"35", x"06", x"76", x"cd", x"e4", x"ad", x"e6",
    x"fd", x"b1", x"05", x"01", x"c9", x"e7", x"14", x"0a",
    x"ee", x"f8", x"f3", x"e4", x"e4", x"2e", x"24", x"0e",
    x"23", x"f1", x"f1", x"14", x"0f", x"9a", x"cd", x"c9",
    x"10", x"09", x"f1", x"f4", x"05", x"fc", x"03", x"f0",
    x"fe", x"c3", x"2c", x"2d", x"1c", x"25", x"19", x"13",
    x"c6", x"07", x"25", x"e8", x"fc", x"38", x"04", x"10",
    x"25", x"04", x"01", x"fc", x"fa", x"fe", x"05", x"04",
    x"01", x"fc", x"1d", x"fd", x"1d", x"27", x"1e", x"02",
    x"fa", x"fa", x"e4", x"1e", x"1e", x"35", x"0a", x"28",
    x"20", x"49", x"1c", x"d4", x"f3", x"00", x"e1", x"e3",
    x"14", x"07", x"c0", x"0d", x"1a", x"dd", x"e2", x"d8",
    x"40", x"ea", x"09", x"00", x"06", x"2a", x"da", x"ee",
    x"f1", x"15", x"11", x"01", x"1b", x"0a", x"0c", x"24",
    x"20", x"33", x"44", x"08", x"f9", x"11", x"e9", x"02",
    x"4e", x"11", x"0a", x"25", x"2c", x"07", x"0a", x"1b",
    x"10", x"ff", x"07", x"f7", x"b2", x"02", x"f7", x"ca",
    x"05", x"28", x"3f", x"0a", x"15", x"48", x"ed", x"0d",
    x"2e", x"f2", x"d5", x"07", x"08", x"f8", x"09", x"08",
    x"12", x"01", x"05", x"04", x"19", x"f1", x"ed", x"25",
    x"ee", x"e7", x"ef", x"07", x"0e", x"b8", x"a7", x"a6",
    x"cf", x"ab", x"c3", x"e1", x"f7", x"00", x"3b", x"56",
    x"39", x"29", x"3b", x"47", x"3e", x"38", x"10", x"11",
    x"0a", x"17", x"05", x"05", x"17", x"e9", x"04", x"1c",
    x"e1", x"08", x"e5", x"cb", x"f2", x"cb", x"a6", x"e0",
    x"e8", x"36", x"35", x"3f", x"19", x"2a", x"55", x"df",
    x"cd", x"a0", x"b1", x"c3", x"aa", x"74", x"a0", x"d0",
    x"3a", x"be", x"ed", x"1f", x"2c", x"28", x"19", x"19",
    x"f5", x"cb", x"14", x"1d", x"fb", x"01", x"09", x"00",
    x"fc", x"f9", x"f8", x"f9", x"00", x"2d", x"2c", x"1e",
    x"0c", x"07", x"2e", x"3f", x"1a", x"18", x"e7", x"03",
    x"34", x"10", x"39", x"1f", x"46", x"25", x"2f", x"24",
    x"0f", x"01", x"09", x"0c", x"05", x"05", x"fb", x"01",
    x"01", x"fb", x"fc", x"ff", x"00", x"03", x"fb", x"00",
    x"fa", x"3e", x"2d", x"37", x"49", x"0b", x"03", x"40",
    x"1c", x"0e", x"38", x"42", x"3e", x"3d", x"34", x"2d",
    x"54", x"21", x"3f", x"10", x"0a", x"f5", x"57", x"02",
    x"10", x"6d", x"29", x"1c", x"fe", x"06", x"dc", x"fd",
    x"f4", x"14", x"f5", x"16", x"19", x"2f", x"25", x"12",
    x"15", x"27", x"58", x"fc", x"06", x"33", x"f7", x"00",
    x"05", x"b5", x"f6", x"16", x"ef", x"e3", x"df", x"fa",
    x"10", x"28", x"1f", x"fe", x"16", x"48", x"16", x"f5",
    x"ff", x"04", x"fe", x"00", x"fe", x"03", x"02", x"03",
    x"f9", x"fe", x"04", x"06", x"04", x"00", x"fe", x"fa",
    x"ff", x"01", x"e3", x"e4", x"0e", x"e3", x"01", x"0c",
    x"05", x"d9", x"0a", x"e5", x"fa", x"aa", x"0a", x"0d",
    x"0b", x"f9", x"f3", x"02", x"d5", x"07", x"13", x"fc",
    x"e5", x"01", x"c2", x"db", x"e1", x"c1", x"ca", x"e2",
    x"e9", x"b0", x"e4", x"f7", x"d8", x"7c", x"0a", x"d7",
    x"99", x"3d", x"04", x"07", x"25", x"fb", x"c8", x"d1",
    x"ac", x"a5", x"aa", x"c3", x"ef", x"01", x"f5", x"22",
    x"d7", x"e7", x"d6", x"b1", x"f2", x"06", x"87", x"3e",
    x"30", x"11", x"0d", x"d5", x"00", x"0b", x"02", x"c5",
    x"ca", x"05", x"ac", x"ef", x"e3", x"20", x"d5", x"c7",
    x"41", x"c5", x"c6", x"1b", x"07", x"06", x"05", x"f9",
    x"06", x"ca", x"c4", x"f4", x"21", x"32", x"3b", x"59",
    x"0c", x"25", x"35", x"06", x"ed", x"d3", x"37", x"1d",
    x"31", x"28", x"25", x"2a", x"01", x"be", x"27", x"20",
    x"2d", x"02", x"0a", x"f3", x"b8", x"f9", x"06", x"d8",
    x"a0", x"ad", x"c1", x"ba", x"a3", x"64", x"aa", x"c8",
    x"fc", x"01", x"fc", x"fc", x"fa", x"01", x"ff", x"fe",
    x"fd", x"ff", x"f9", x"00", x"01", x"01", x"fb", x"02",
    x"01", x"fb", x"fb", x"02", x"fc", x"fd", x"fe", x"f8",
    x"03", x"fd", x"fc", x"f6", x"fc", x"fd", x"fc", x"f9",
    x"fb", x"fc", x"fd", x"fb", x"fe", x"fb", x"f9", x"03",
    x"00", x"02", x"02", x"04", x"fc", x"00", x"f7", x"fc",
    x"04", x"fd", x"fe", x"fb", x"fc", x"fb", x"fb", x"ff",
    x"fb", x"fd", x"03", x"fb", x"fb", x"ff", x"02", x"fd",
    x"03", x"01", x"00", x"00", x"00", x"fc", x"f7", x"04",
    x"00", x"fd", x"ff", x"00", x"f7", x"f9", x"02", x"fa",
    x"fa", x"fb", x"f9", x"f6", x"fe", x"fc", x"fe", x"04",
    x"01", x"fc", x"fb", x"ff", x"02", x"03", x"fc", x"03",
    x"00", x"ff", x"ff", x"01", x"fd", x"fa", x"04", x"fd",
    x"01", x"01", x"04", x"fe", x"fd", x"00", x"fe", x"02",
    x"f9", x"f7", x"fe", x"fb", x"ff", x"fe", x"fd", x"fe",
    x"f9", x"f6", x"01", x"04", x"00", x"fb", x"fb", x"f8",
    x"00", x"fb", x"f9", x"02", x"fb", x"02", x"fb", x"fb",
    x"01", x"fb", x"fe", x"ff", x"02", x"fd", x"fd", x"01",
    x"fd", x"ff", x"00", x"fb", x"fc", x"00", x"01", x"ff",
    x"fe", x"00", x"02", x"03", x"fb", x"01", x"fc", x"fd",
    x"01", x"02", x"00", x"03", x"fa", x"fc", x"f6", x"02",
    x"ff", x"fa", x"04", x"fd", x"fa", x"00", x"01", x"ff",
    x"fc", x"fd", x"fd", x"00", x"fd", x"ff", x"01", x"fd",
    x"fc", x"fe", x"03", x"fe", x"ff", x"f7", x"fd", x"03",
    x"04", x"02", x"00", x"fd", x"fb", x"fd", x"fd", x"03",
    x"fc", x"00", x"fc", x"fc", x"fd", x"fd", x"01", x"f7",
    x"ff", x"ff", x"00", x"04", x"fb", x"03", x"fd", x"fb",
    x"04", x"00", x"fa", x"fd", x"02", x"fc", x"00", x"02",
    x"fd", x"00", x"f7", x"02", x"fb", x"fd", x"fe", x"fd",
    x"fd", x"02", x"fd", x"01", x"fa", x"00", x"02", x"fa",
    x"fa", x"03", x"fa", x"ff", x"02", x"01", x"ff", x"05",
    x"03", x"02", x"03", x"03", x"f6", x"f8", x"04", x"fd",
    x"03", x"04", x"fb", x"fa", x"04", x"fe", x"f9", x"fe",
    x"04", x"01", x"00", x"01", x"fd", x"02", x"fb", x"fb",
    x"fb", x"00", x"03", x"03", x"fb", x"fd", x"f6", x"fa",
    x"fd", x"02", x"fd", x"01", x"f9", x"01", x"ff", x"01",
    x"00", x"03", x"03", x"fb", x"fb", x"01", x"fe", x"f6",
    x"ff", x"00", x"fd", x"fa", x"05", x"fd", x"fb", x"04",
    x"fe", x"fb", x"f7", x"00", x"03", x"f9", x"ff", x"00",
    x"02", x"fe", x"fe", x"fa", x"00", x"fe", x"03", x"00",
    x"01", x"fa", x"ff", x"02", x"02", x"03", x"02", x"01",
    x"fe", x"00", x"00", x"02", x"00", x"fc", x"fa", x"01",
    x"fd", x"00", x"fd", x"02", x"fe", x"fb", x"fd", x"fb",
    x"fb", x"fa", x"00", x"03", x"ff", x"fe", x"00", x"fa",
    x"ff", x"fa", x"f6", x"00", x"01", x"fe", x"ff", x"fe",
    x"fe", x"03", x"fe", x"01", x"01", x"fc", x"ff", x"fc",
    x"04", x"ff", x"01", x"fe", x"fd", x"00", x"fc", x"ff",
    x"fe", x"fe", x"04", x"fc", x"02", x"fd", x"fd", x"f9",
    x"fb", x"fb", x"fe", x"fa", x"f6", x"ff", x"02", x"fb",
    x"fd", x"fd", x"01", x"01", x"fc", x"fe", x"00", x"fb",
    x"fa", x"fc", x"fd", x"01", x"fd", x"f8", x"fa", x"fe",
    x"f8", x"ff", x"fc", x"02", x"00", x"fc", x"fc", x"fc",
    x"ff", x"00", x"f9", x"ff", x"01", x"fd", x"01", x"f9",
    x"f8", x"04", x"fc", x"00", x"fe", x"fe", x"ff", x"fd",
    x"05", x"03", x"fb", x"00", x"02", x"fe", x"04", x"04",
    x"04", x"fe", x"00", x"02", x"03", x"fb", x"02", x"fe",
    x"fb", x"02", x"f6", x"fc", x"04", x"fb", x"fe", x"fe",
    x"ff", x"fa", x"fd", x"fe", x"fe", x"fe", x"fb", x"ff",
    x"fa", x"04", x"f9", x"ff", x"f9", x"fe", x"fd", x"03",
    x"fa", x"fd", x"03", x"04", x"fb", x"fb", x"fb", x"ff",
    x"fb", x"f8", x"fd", x"fe", x"00", x"fd", x"01", x"ff",
    x"03", x"00", x"00", x"fd", x"03", x"fd", x"fc", x"01",
    x"fb", x"fe", x"f6", x"ff", x"02", x"fb", x"02", x"fa",
    x"01", x"fd", x"02", x"03", x"fe", x"fb", x"fa", x"01",
    x"fb", x"fa", x"04", x"fa", x"00", x"ff", x"fa", x"fa",
    x"fd", x"fc", x"fb", x"00", x"fe", x"f8", x"02", x"00",
    x"00", x"fd", x"ff", x"fc", x"f9", x"00", x"fd", x"fc",
    x"fb", x"04", x"fc", x"fd", x"ff", x"fb", x"fb", x"fe",
    x"01", x"ff", x"fb", x"fd", x"00", x"fc", x"fb", x"00",
    x"fc", x"02", x"ff", x"fb", x"fe", x"ff", x"fd", x"fb",
    x"02", x"fc", x"fd", x"fa", x"fc", x"fe", x"fc", x"f7",
    x"fa", x"00", x"f8", x"ff", x"fa", x"fc", x"fa", x"fd",
    x"27", x"11", x"4c", x"06", x"08", x"f3", x"d1", x"f8",
    x"08", x"59", x"1f", x"31", x"f0", x"22", x"2d", x"ed",
    x"f4", x"31", x"32", x"21", x"2a", x"26", x"00", x"11",
    x"1c", x"0d", x"34", x"d8", x"b3", x"ca", x"f7", x"f9",
    x"b7", x"e6", x"e6", x"b1", x"1d", x"f4", x"16", x"35",
    x"34", x"53", x"4a", x"4c", x"67", x"ea", x"cb", x"00",
    x"e5", x"d9", x"00", x"d8", x"e6", x"df", x"11", x"e9",
    x"0f", x"dc", x"c6", x"03", x"88", x"d8", x"e5", x"14",
    x"0c", x"35", x"fa", x"0e", x"1e", x"f2", x"05", x"1b",
    x"26", x"38", x"64", x"1d", x"1b", x"2d", x"0e", x"1a",
    x"40", x"11", x"fd", x"fb", x"35", x"15", x"b4", x"13",
    x"d1", x"a6", x"e3", x"fc", x"df", x"a6", x"e5", x"d5",
    x"27", x"57", x"33", x"00", x"c4", x"e6", x"fd", x"be",
    x"c7", x"07", x"da", x"b8", x"0e", x"34", x"3b", x"ed",
    x"2f", x"41", x"15", x"14", x"34", x"34", x"2d", x"4d",
    x"23", x"27", x"11", x"ce", x"f8", x"41", x"e8", x"d9",
    x"e6", x"0b", x"d2", x"e8", x"28", x"f4", x"ce", x"20",
    x"f7", x"d5", x"1f", x"e0", x"d5", x"24", x"d8", x"81",
    x"c8", x"f0", x"e4", x"f9", x"e6", x"bd", x"00", x"fe",
    x"f0", x"01", x"04", x"ff", x"fe", x"fc", x"fd", x"02",
    x"fb", x"03", x"f1", x"30", x"d8", x"ce", x"c4", x"ef",
    x"e3", x"ea", x"0a", x"e3", x"1d", x"09", x"f9", x"1d",
    x"fa", x"c4", x"e7", x"17", x"15", x"3e", x"33", x"f7",
    x"17", x"49", x"ef", x"eb", x"4b", x"07", x"04", x"f5",
    x"0b", x"03", x"10", x"52", x"40", x"66", x"fa", x"e7",
    x"03", x"d5", x"c6", x"ca", x"cb", x"ab", x"29", x"47",
    x"f9", x"ed", x"3e", x"32", x"1a", x"f3", x"1d", x"4e",
    x"f4", x"3c", x"41", x"ae", x"12", x"35", x"08", x"9c",
    x"e0", x"0c", x"09", x"fb", x"a5", x"eb", x"f3", x"e4",
    x"e9", x"1b", x"22", x"11", x"0c", x"0b", x"0a", x"1a",
    x"3e", x"2b", x"6b", x"08", x"01", x"02", x"fe", x"fc",
    x"07", x"03", x"fd", x"0d", x"07", x"d1", x"e8", x"16",
    x"01", x"f7", x"04", x"1c", x"0e", x"09", x"f5", x"d8",
    x"f3", x"15", x"f6", x"f7", x"f0", x"d3", x"30", x"1a",
    x"2b", x"1c", x"29", x"18", x"05", x"14", x"28", x"02",
    x"f9", x"fe", x"ed", x"0f", x"08", x"14", x"e4", x"ef",
    x"20", x"e8", x"c1", x"ca", x"b5", x"d8", x"f0", x"e6",
    x"c2", x"05", x"06", x"f8", x"3e", x"11", x"ed", x"00",
    x"f2", x"0f", x"17", x"15", x"01", x"00", x"11", x"11",
    x"00", x"0f", x"0f", x"03", x"28", x"16", x"fd", x"3a",
    x"01", x"c5", x"7d", x"2b", x"05", x"03", x"fb", x"ff",
    x"0e", x"0a", x"06", x"08", x"02", x"3e", x"15", x"01",
    x"22", x"20", x"10", x"0c", x"1e", x"00", x"e0", x"f2",
    x"05", x"3d", x"d8", x"aa", x"e6", x"7a", x"8f", x"f4",
    x"eb", x"1a", x"c6", x"ab", x"b8", x"e5", x"9a", x"8e",
    x"ff", x"03", x"06", x"fd", x"02", x"fe", x"ff", x"04",
    x"fb", x"3e", x"28", x"41", x"17", x"17", x"31", x"2d",
    x"2a", x"0b", x"29", x"09", x"10", x"33", x"0c", x"24",
    x"5b", x"1c", x"19", x"22", x"21", x"17", x"49", x"3e",
    x"22", x"00", x"3e", x"35", x"55", x"47", x"3f", x"13",
    x"0e", x"0a", x"00", x"0f", x"1e", x"20", x"25", x"50",
    x"15", x"0e", x"16", x"27", x"0e", x"02", x"30", x"1a",
    x"53", x"2c", x"d7", x"c4", x"08", x"f0", x"ce", x"29",
    x"f1", x"ea", x"03", x"e0", x"e0", x"f1", x"f5", x"ed",
    x"02", x"fa", x"01", x"fd", x"fe", x"ff", x"fc", x"05",
    x"fd", x"01", x"03", x"fd", x"01", x"fb", x"04", x"04",
    x"06", x"ff", x"ce", x"d4", x"d3", x"f0", x"e5", x"d5",
    x"1b", x"07", x"f7", x"e9", x"b4", x"be", x"d3", x"bc",
    x"b9", x"d4", x"f8", x"d1", x"17", x"00", x"ec", x"10",
    x"07", x"f7", x"c5", x"cc", x"f4", x"f5", x"f1", x"fb",
    x"0a", x"07", x"01", x"08", x"1a", x"43", x"fe", x"e5",
    x"ed", x"f1", x"e9", x"10", x"fa", x"fb", x"dd", x"5d",
    x"12", x"0a", x"dc", x"e9", x"0a", x"92", x"c6", x"c2",
    x"f2", x"1c", x"f8", x"f7", x"cd", x"d1", x"ed", x"02",
    x"01", x"07", x"00", x"08", x"34", x"0a", x"3b", x"e8",
    x"e8", x"54", x"e2", x"e9", x"17", x"cf", x"ac", x"dd",
    x"e1", x"bd", x"ac", x"f0", x"d1", x"e4", x"22", x"1f",
    x"34", x"f5", x"27", x"20", x"11", x"16", x"32", x"36",
    x"fd", x"09", x"20", x"fc", x"14", x"18", x"1b", x"04",
    x"ed", x"11", x"ec", x"44", x"18", x"1b", x"0d", x"32",
    x"23", x"0d", x"23", x"39", x"0a", x"17", x"49", x"13",
    x"fd", x"2c", x"e1", x"f3", x"08", x"cc", x"da", x"f3",
    x"ec", x"2b", x"52", x"0b", x"0e", x"0e", x"06", x"db",
    x"23", x"3f", x"2e", x"38", x"d5", x"11", x"1c", x"09",
    x"3e", x"1d", x"fb", x"01", x"0d", x"0a", x"2a", x"1c",
    x"3c", x"31", x"f2", x"8c", x"2e", x"cd", x"b1", x"cc",
    x"dc", x"da", x"be", x"c5", x"f2", x"10", x"ef", x"29",
    x"4d", x"5b", x"23", x"e8", x"31", x"e1", x"e9", x"06",
    x"93", x"02", x"3f", x"b3", x"1d", x"11", x"08", x"4e",
    x"2d", x"c2", x"a8", x"cc", x"73", x"5e", x"19", x"2f",
    x"1c", x"24", x"0a", x"02", x"26", x"1c", x"0d", x"0b",
    x"21", x"33", x"64", x"f1", x"0d", x"52", x"13", x"2a",
    x"4d", x"12", x"dd", x"b7", x"de", x"c6", x"9c", x"9f",
    x"b1", x"a6", x"2c", x"28", x"f2", x"bd", x"ec", x"f9",
    x"e4", x"2a", x"0f", x"53", x"1f", x"fa", x"39", x"00",
    x"ef", x"4c", x"d2", x"c0", x"3a", x"12", x"1a", x"27",
    x"0f", x"fb", x"0d", x"24", x"23", x"2a", x"4b", x"29",
    x"0c", x"de", x"8d", x"f1", x"c7", x"eb", x"c4", x"df",
    x"14", x"1a", x"fa", x"19", x"23", x"28", x"06", x"47",
    x"31", x"ee", x"42", x"49", x"c0", x"3b", x"db", x"8b",
    x"24", x"07", x"f7", x"35", x"e0", x"dc", x"2c", x"f2",
    x"4e", x"04", x"00", x"04", x"fc", x"03", x"04", x"fb",
    x"01", x"01", x"d9", x"ed", x"09", x"fc", x"cd", x"ed",
    x"fc", x"f8", x"0a", x"07", x"2a", x"2e", x"e8", x"04",
    x"20", x"a7", x"9e", x"f6", x"47", x"87", x"00", x"0a",
    x"d0", x"fa", x"15", x"fa", x"17", x"21", x"2b", x"11",
    x"30", x"11", x"0a", x"4f", x"fb", x"46", x"f5", x"10",
    x"2c", x"ef", x"0c", x"f5", x"3e", x"2b", x"1b", x"1e",
    x"1e", x"2d", x"2d", x"3b", x"3a", x"54", x"15", x"1c",
    x"d7", x"62", x"23", x"ed", x"15", x"fe", x"ec", x"eb",
    x"fc", x"30", x"17", x"eb", x"b9", x"d9", x"bd", x"d7",
    x"ea", x"f8", x"e2", x"f5", x"16", x"0b", x"18", x"2d",
    x"2d", x"0b", x"6a", x"04", x"09", x"03", x"fa", x"02",
    x"02", x"fb", x"03", x"07", x"05", x"11", x"0d", x"10",
    x"10", x"17", x"06", x"0f", x"28", x"15", x"01", x"f3",
    x"f4", x"f8", x"ed", x"18", x"b9", x"d1", x"ce", x"d2",
    x"fc", x"eb", x"da", x"ed", x"f1", x"ef", x"00", x"2d",
    x"3e", x"10", x"03", x"13", x"23", x"f1", x"f2", x"e9",
    x"34", x"30", x"1c", x"dd", x"da", x"da", x"f4", x"f1",
    x"eb", x"29", x"d9", x"c1", x"d7", x"a7", x"ba", x"d9",
    x"dc", x"2c", x"29", x"4f", x"4a", x"13", x"36", x"33",
    x"0d", x"24", x"2d", x"f7", x"38", x"f6", x"e0", x"df",
    x"da", x"de", x"ff", x"01", x"05", x"09", x"03", x"03",
    x"05", x"0b", x"08", x"09", x"07", x"45", x"f8", x"d8",
    x"30", x"c0", x"d0", x"ee", x"e9", x"ca", x"d3", x"f6",
    x"01", x"15", x"20", x"fd", x"4c", x"f0", x"da", x"22",
    x"4f", x"f2", x"06", x"c9", x"dc", x"da", x"ed", x"b4",
    x"fc", x"fe", x"03", x"fd", x"03", x"02", x"02", x"01",
    x"fc", x"da", x"d2", x"ee", x"e7", x"d9", x"fd", x"1d",
    x"cc", x"ec", x"0e", x"07", x"01", x"00", x"08", x"15",
    x"19", x"0a", x"f6", x"2a", x"fb", x"16", x"0e", x"0e",
    x"25", x"05", x"19", x"32", x"59", x"1d", x"0f", x"74",
    x"32", x"01", x"45", x"45", x"2b", x"e8", x"1c", x"20",
    x"11", x"fd", x"f0", x"16", x"fe", x"fe", x"1d", x"43",
    x"3f", x"e2", x"fd", x"1d", x"f8", x"e8", x"fb", x"23",
    x"2a", x"32", x"24", x"30", x"4e", x"33", x"20", x"2a",
    x"03", x"fd", x"03", x"03", x"fe", x"02", x"fd", x"04",
    x"fa", x"fe", x"ff", x"02", x"02", x"fd", x"01", x"01",
    x"02", x"f9", x"ff", x"e4", x"00", x"1c", x"1b", x"32",
    x"52", x"2d", x"42", x"e2", x"d7", x"12", x"ee", x"e4",
    x"bd", x"f3", x"e8", x"ca", x"d2", x"dd", x"e7", x"c3",
    x"a6", x"eb", x"bd", x"9f", x"ea", x"ec", x"ff", x"ef",
    x"44", x"2f", x"12", x"5e", x"3f", x"19", x"f9", x"2b",
    x"f2", x"0e", x"03", x"04", x"04", x"fb", x"23", x"1d",
    x"1b", x"1e", x"cb", x"d3", x"e0", x"b3", x"bc", x"b4",
    x"dc", x"0a", x"30", x"d1", x"c1", x"e7", x"43", x"bc",
    x"ec", x"f4", x"0d", x"ed", x"de", x"fe", x"38", x"ed",
    x"1c", x"26", x"f6", x"e6", x"f6", x"eb", x"b1", x"e5",
    x"01", x"c0", x"c8", x"ff", x"f7", x"f8", x"0e", x"1f",
    x"0e", x"f5", x"2d", x"27", x"30", x"e6", x"f2", x"04",
    x"fd", x"01", x"f0", x"ed", x"05", x"0e", x"11", x"fb",
    x"f1", x"14", x"02", x"ed", x"17", x"14", x"1d", x"04",
    x"07", x"21", x"04", x"11", x"51", x"fc", x"ee", x"11",
    x"0c", x"22", x"27", x"10", x"17", x"19", x"2f", x"59",
    x"08", x"0d", x"85", x"f0", x"f3", x"0f", x"16", x"c9",
    x"7b", x"1d", x"f3", x"fb", x"19", x"09", x"ea", x"3d",
    x"31", x"14", x"22", x"20", x"f5", x"17", x"09", x"14",
    x"1d", x"1b", x"3e", x"0b", x"da", x"cf", x"d9", x"ce",
    x"fa", x"9f", x"b9", x"ee", x"b7", x"cf", x"c8", x"fc",
    x"10", x"ed", x"05", x"11", x"fe", x"e9", x"1f", x"2d",
    x"c5", x"0c", x"5a", x"ff", x"35", x"4a", x"f8", x"ed",
    x"f6", x"27", x"ef", x"eb", x"de", x"85", x"ba", x"da",
    x"dc", x"61", x"04", x"0e", x"01", x"0d", x"07", x"cc",
    x"db", x"a3", x"b1", x"c3", x"ca", x"c7", x"d2", x"f8",
    x"d1", x"e8", x"e4", x"f3", x"03", x"0c", x"32", x"27",
    x"17", x"65", x"02", x"f8", x"15", x"a8", x"c8", x"15",
    x"20", x"2b", x"fd", x"14", x"20", x"19", x"1d", x"15",
    x"24", x"72", x"db", x"da", x"ff", x"db", x"b8", x"02",
    x"0b", x"e2", x"38", x"f8", x"22", x"de", x"16", x"85",
    x"17", x"28", x"1f", x"35", x"11", x"01", x"23", x"13",
    x"d7", x"f8", x"10", x"ed", x"05", x"11", x"10", x"54",
    x"1f", x"f7", x"01", x"2d", x"57", x"16", x"31", x"40",
    x"38", x"1b", x"34", x"56", x"29", x"20", x"1f", x"2e",
    x"ff", x"04", x"00", x"05", x"01", x"fe", x"04", x"fe",
    x"fd", x"05", x"d2", x"14", x"38", x"09", x"2d", x"31",
    x"28", x"39", x"17", x"c0", x"f1", x"04", x"dd", x"f1",
    x"f9", x"15", x"ff", x"ed", x"d6", x"03", x"30", x"ff",
    x"00", x"12", x"f9", x"30", x"04", x"de", x"ef", x"e7",
    x"fb", x"f6", x"e9", x"59", x"11", x"dd", x"27", x"42",
    x"5b", x"1d", x"48", x"2b", x"33", x"45", x"e7", x"a0",
    x"20", x"13", x"a2", x"02", x"1a", x"fb", x"0a", x"d3",
    x"15", x"fe", x"11", x"26", x"f8", x"ee", x"b7", x"f9",
    x"f1", x"2f", x"30", x"0c", x"63", x"32", x"08", x"3b",
    x"29", x"e9", x"ca", x"cd", x"de", x"c8", x"c6", x"91",
    x"8f", x"35", x"b2", x"05", x"0a", x"03", x"fd", x"fd",
    x"03", x"01", x"01", x"04", x"d6", x"ea", x"c7", x"f5",
    x"e9", x"f1", x"0b", x"fb", x"0d", x"2a", x"12", x"04",
    x"2d", x"fa", x"cb", x"05", x"de", x"bf", x"e0", x"05",
    x"fd", x"fc", x"d6", x"e5", x"0d", x"05", x"03", x"ce",
    x"e2", x"dc", x"e4", x"16", x"1a", x"0b", x"0a", x"13",
    x"d4", x"15", x"28", x"00", x"ed", x"05", x"eb", x"f7",
    x"fb", x"d4", x"e1", x"02", x"fc", x"f7", x"f3", x"32",
    x"f7", x"e5", x"39", x"45", x"82", x"01", x"1e", x"46",
    x"f1", x"2a", x"20", x"f8", x"f9", x"d8", x"d7", x"c6",
    x"f4", x"1d", x"e0", x"c9", x"f9", x"f9", x"04", x"f9",
    x"f6", x"f9", x"fb", x"f8", x"f5", x"17", x"fd", x"07",
    x"44", x"f6", x"13", x"28", x"13", x"e7", x"27", x"17",
    x"32", x"61", x"0d", x"0d", x"39", x"fa", x"0b", x"14",
    x"bf", x"e2", x"fa", x"1c", x"00", x"2b", x"fb", x"03",
    x"fe", x"fe", x"04", x"fc", x"fc", x"01", x"fe", x"02",
    x"04", x"3c", x"b1", x"a5", x"45", x"bd", x"b8", x"2b",
    x"0e", x"dd", x"1c", x"e9", x"0b", x"01", x"00", x"fc",
    x"08", x"e9", x"d2", x"1e", x"04", x"e9", x"2f", x"ce",
    x"cb", x"24", x"e1", x"c5", x"36", x"43", x"5d", x"1c",
    x"20", x"25", x"51", x"35", x"4f", x"dc", x"d1", x"cd",
    x"cb", x"94", x"b1", x"f8", x"c4", x"c2", x"c2", x"f4",
    x"70", x"3a", x"01", x"f1", x"2f", x"27", x"1a", x"df",
    x"13", x"ff", x"03", x"16", x"14", x"fe", x"17", x"03",
    x"01", x"03", x"fe", x"02", x"06", x"00", x"08", x"fa",
    x"04", x"fe", x"05", x"03", x"01", x"fd", x"fd", x"08",
    x"00", x"09", x"1b", x"29", x"00", x"e8", x"f9", x"01",
    x"e1", x"e9", x"0c", x"e5", x"fd", x"0c", x"d5", x"ee",
    x"01", x"d0", x"c0", x"da", x"c9", x"d0", x"00", x"db",
    x"ca", x"df", x"f6", x"f6", x"e2", x"20", x"1f", x"fb",
    x"1a", x"16", x"09", x"78", x"57", x"ea", x"2f", x"03",
    x"11", x"e6", x"06", x"05", x"0e", x"0a", x"e7", x"bc",
    x"d8", x"03", x"d4", x"96", x"ce", x"b3", x"ae", x"b9",
    x"02", x"17", x"37", x"f3", x"18", x"14", x"53", x"05",
    x"25", x"36", x"ff", x"cf", x"1c", x"e4", x"ea", x"1c",
    x"e1", x"10", x"26", x"0d", x"01", x"10", x"1b", x"17",
    x"e3", x"3a", x"25", x"38", x"05", x"fc", x"40", x"19",
    x"33", x"8f", x"6f", x"55", x"11", x"80", x"17", x"da",
    x"34", x"3c", x"14", x"1b", x"0c", x"e4", x"fc", x"2c",
    x"f8", x"e5", x"dc", x"07", x"20", x"00", x"30", x"0d",
    x"f6", x"15", x"fc", x"f8", x"00", x"03", x"dd", x"0c",
    x"2b", x"24", x"e2", x"00", x"2b", x"1d", x"52", x"51",
    x"00", x"09", x"3d", x"f2", x"ea", x"de", x"0b", x"3e",
    x"46", x"25", x"f5", x"12", x"e1", x"02", x"09", x"07",
    x"20", x"ff", x"d0", x"23", x"21", x"3d", x"1d", x"e5",
    x"01", x"e4", x"be", x"16", x"fb", x"c7", x"0b", x"e8",
    x"ee", x"f4", x"f4", x"cb", x"c5", x"de", x"cd", x"20",
    x"08", x"f1", x"13", x"d8", x"fa", x"ff", x"d5", x"ec",
    x"1a", x"19", x"f6", x"8a", x"fa", x"b7", x"61", x"38",
    x"4f", x"e2", x"0d", x"13", x"35", x"23", x"00", x"de",
    x"fb", x"3e", x"66", x"61", x"c0", x"be", x"ca", x"13",
    x"f4", x"e4", x"f5", x"91", x"8f", x"87", x"0c", x"02",
    x"3b", x"dc", x"05", x"e8", x"ca", x"d7", x"cb", x"bd",
    x"9b", x"0d", x"2e", x"47", x"4c", x"f2", x"40", x"25",
    x"34", x"01", x"fe", x"16", x"f1", x"1e", x"fd", x"fb",
    x"2b", x"1b", x"02", x"2b", x"23", x"b4", x"c3", x"08",
    x"1d", x"25", x"3a", x"33", x"03", x"01", x"00", x"1f",
    x"e7", x"c6", x"24", x"fc", x"f6", x"11", x"ef", x"19",
    x"f4", x"18", x"09", x"da", x"c3", x"d3", x"d3", x"1b",
    x"f8", x"fd", x"e4", x"d3", x"19", x"c5", x"f5", x"fa",
    x"d6", x"f4", x"fe", x"e0", x"eb", x"f2", x"0b", x"07",
    x"f8", x"ff", x"01", x"ff", x"fe", x"01", x"05", x"00",
    x"ff", x"01", x"db", x"e6", x"d4", x"cc", x"04", x"06",
    x"42", x"d3", x"e4", x"0d", x"1e", x"e6", x"27", x"04",
    x"e4", x"e7", x"18", x"29", x"d8", x"ed", x"f4", x"ca",
    x"05", x"f8", x"02", x"15", x"f9", x"b7", x"f2", x"f2",
    x"29", x"1c", x"39", x"d8", x"02", x"e2", x"d9", x"0f",
    x"1f", x"de", x"fe", x"fd", x"f8", x"0c", x"12", x"f9",
    x"90", x"0d", x"23", x"00", x"fe", x"0e", x"e4", x"11",
    x"e9", x"de", x"2d", x"ba", x"17", x"14", x"3c", x"f9",
    x"fa", x"cb", x"ff", x"f9", x"b3", x"f7", x"10", x"1e",
    x"3c", x"0a", x"ce", x"14", x"e0", x"c8", x"1a", x"2c",
    x"17", x"32", x"3b", x"f8", x"fc", x"fa", x"f7", x"f9",
    x"fd", x"fa", x"fc", x"ff", x"ed", x"e6", x"dd", x"bf",
    x"ae", x"df", x"d5", x"be", x"e5", x"de", x"d4", x"39",
    x"03", x"14", x"26", x"57", x"0a", x"44", x"df", x"d8",
    x"ce", x"07", x"04", x"d7", x"c8", x"8c", x"ca", x"b5",
    x"a4", x"c2", x"ca", x"d6", x"ed", x"fb", x"f0", x"fb",
    x"b3", x"cc", x"11", x"e0", x"f6", x"3f", x"3f", x"2c",
    x"fd", x"f2", x"12", x"09", x"b4", x"e5", x"e9", x"d6",
    x"b5", x"19", x"9b", x"fa", x"44", x"fc", x"21", x"07",
    x"16", x"06", x"e9", x"e2", x"f2", x"00", x"f4", x"ca",
    x"a3", x"e7", x"0c", x"18", x"03", x"ff", x"01", x"09",
    x"03", x"fe", x"08", x"04", x"0f", x"fe", x"de", x"f5",
    x"e6", x"10", x"2b", x"cf", x"2a", x"30", x"f7", x"0d",
    x"1a", x"08", x"e6", x"cb", x"26", x"f1", x"ed", x"c3",
    x"14", x"1b", x"cc", x"1a", x"03", x"45", x"29", x"24",
    x"02", x"00", x"00", x"05", x"fe", x"00", x"01", x"02",
    x"00", x"01", x"f0", x"ec", x"0f", x"ed", x"d7", x"c5",
    x"fc", x"12", x"23", x"f0", x"d9", x"29", x"05", x"f4",
    x"29", x"26", x"3f", x"23", x"36", x"26", x"c0", x"fb",
    x"ff", x"08", x"26", x"09", x"e6", x"c7", x"d1", x"e3",
    x"e8", x"2e", x"12", x"1a", x"2e", x"e7", x"f5", x"22",
    x"30", x"52", x"3e", x"21", x"1e", x"24", x"a6", x"03",
    x"5c", x"aa", x"2d", x"fc", x"93", x"f7", x"f5", x"11",
    x"d8", x"f6", x"23", x"06", x"37", x"d8", x"1f", x"fe",
    x"fd", x"03", x"00", x"03", x"05", x"04", x"05", x"02",
    x"fb", x"05", x"00", x"fc", x"00", x"ff", x"fb", x"ff",
    x"fe", x"03", x"d8", x"f3", x"f3", x"fd", x"2d", x"19",
    x"33", x"41", x"1a", x"f1", x"10", x"05", x"4d", x"3d",
    x"00", x"2d", x"f1", x"a7", x"fe", x"10", x"01", x"0a",
    x"fc", x"0f", x"02", x"bd", x"c3", x"dc", x"dd", x"d5",
    x"db", x"e2", x"da", x"2d", x"f9", x"03", x"c3", x"30",
    x"13", x"dd", x"e9", x"25", x"ae", x"04", x"d7", x"b8",
    x"29", x"4a", x"1c", x"33", x"16", x"6b", x"17", x"3f",
    x"62", x"24", x"05", x"1e", x"0b", x"e4", x"2a", x"22",
    x"ff", x"ba", x"cc", x"db", x"7c", x"2a", x"14", x"fb",
    x"09", x"18", x"21", x"31", x"25", x"30", x"fc", x"17",
    x"1a", x"1b", x"32", x"ea", x"01", x"e6", x"03", x"13",
    x"05", x"fe", x"fb", x"b9", x"03", x"fc", x"a1", x"ec",
    x"50", x"67", x"ec", x"27", x"30", x"d3", x"f8", x"fa",
    x"10", x"09", x"e2", x"f6", x"1d", x"25", x"3c", x"e8",
    x"11", x"db", x"e6", x"f5", x"f8", x"01", x"0b", x"a8",
    x"04", x"2b", x"10", x"4a", x"3d", x"27", x"14", x"ed",
    x"f9", x"1a", x"2a", x"c8", x"03", x"d8", x"aa", x"e8",
    x"59", x"3c", x"05", x"f3", x"05", x"33", x"25", x"04",
    x"0d", x"56", x"27", x"03", x"f9", x"1c", x"0c", x"01",
    x"49", x"20", x"ef", x"06", x"f1", x"e5", x"e5", x"f0",
    x"df", x"8e", x"b0", x"d8", x"e4", x"de", x"da", x"f8",
    x"e1", x"d9", x"c4", x"d2", x"f6", x"00", x"16", x"0b",
    x"ec", x"15", x"25", x"11", x"20", x"3f", x"d8", x"e3",
    x"fe", x"db", x"da", x"ff", x"ca", x"d4", x"de", x"d9",
    x"f0", x"3e", x"d2", x"e7", x"51", x"d2", x"f4", x"30",
    x"d8", x"f3", x"56", x"e9", x"01", x"2f", x"e6", x"05",
    x"40", x"0d", x"0d", x"24", x"45", x"24", x"0f", x"80",
    x"39", x"fb", x"0f", x"e1", x"cd", x"f7", x"c9", x"e1",
    x"5f", x"00", x"26", x"fa", x"2e", x"1b", x"2d", x"27",
    x"08", x"47", x"1a", x"0b", x"a0", x"ef", x"17", x"cc",
    x"1a", x"15", x"e2", x"e2", x"05", x"27", x"2a", x"4f",
    x"19", x"06", x"e7", x"dc", x"fe", x"3c", x"0d", x"f8",
    x"de", x"d9", x"c7", x"d6", x"e2", x"b4", x"c9", x"04",
    x"f0", x"f4", x"d2", x"ed", x"19", x"0f", x"18", x"ff",
    x"a5", x"de", x"f9", x"d7", x"e6", x"13", x"07", x"05",
    x"0d", x"05", x"03", x"02", x"03", x"03", x"03", x"01",
    x"00", x"05", x"da", x"1c", x"21", x"f7", x"17", x"19",
    x"27", x"08", x"2f", x"e6", x"f5", x"f8", x"ee", x"06",
    x"39", x"22", x"2b", x"53", x"1c", x"1d", x"eb", x"d9",
    x"20", x"27", x"ec", x"d4", x"45", x"e2", x"da", x"d8",
    x"22", x"09", x"ec", x"49", x"03", x"2d", x"08", x"01",
    x"03", x"e8", x"f9", x"26", x"a7", x"b2", x"20", x"1a",
    x"d4", x"c5", x"27", x"f1", x"fc", x"bd", x"d8", x"00",
    x"23", x"5b", x"45", x"cc", x"42", x"26", x"fa", x"c5",
    x"f4", x"0e", x"18", x"d8", x"f9", x"0c", x"f9", x"ec",
    x"e0", x"30", x"e9", x"14", x"03", x"cb", x"fa", x"1b",
    x"33", x"2e", x"55", x"06", x"09", x"03", x"07", x"10",
    x"0f", x"0a", x"05", x"f9", x"dc", x"cd", x"d4", x"f6",
    x"be", x"e2", x"ea", x"e4", x"db", x"de", x"c8", x"fd",
    x"e0", x"be", x"e8", x"e7", x"e2", x"f7", x"12", x"4b",
    x"46", x"37", x"4a", x"2a", x"09", x"31", x"1d", x"96",
    x"ca", x"c0", x"ca", x"d7", x"df", x"0f", x"00", x"f4",
    x"0b", x"f5", x"31", x"c2", x"d4", x"c9", x"e0", x"b9",
    x"b6", x"01", x"f3", x"f7", x"0e", x"f2", x"db", x"3b",
    x"1d", x"1e", x"9b", x"f1", x"fe", x"d4", x"e1", x"e1",
    x"b9", x"d3", x"18", x"cd", x"2c", x"1b", x"0b", x"0e",
    x"17", x"d9", x"07", x"ed", x"f6", x"06", x"0a", x"f5",
    x"09", x"07", x"00", x"ff", x"06", x"35", x"00", x"f0",
    x"e4", x"fe", x"fd", x"e5", x"06", x"ee", x"e6", x"f0",
    x"fa", x"dc", x"d7", x"ea", x"cc", x"e5", x"c0", x"da",
    x"e2", x"f5", x"c5", x"d9", x"07", x"6f", x"8d", x"bc",
    x"fc", x"fc", x"01", x"ff", x"ff", x"02", x"00", x"02",
    x"fb", x"6d", x"ff", x"fc", x"2f", x"15", x"01", x"48",
    x"17", x"38", x"1e", x"32", x"0c", x"4a", x"40", x"21",
    x"3a", x"e4", x"30", x"41", x"10", x"07", x"3d", x"33",
    x"25", x"6d", x"45", x"29", x"e8", x"fe", x"1f", x"14",
    x"05", x"18", x"ef", x"f0", x"ec", x"b3", x"f5", x"2b",
    x"f1", x"f4", x"fe", x"01", x"09", x"14", x"d0", x"00",
    x"02", x"ff", x"ce", x"d5", x"21", x"f4", x"ef", x"4a",
    x"06", x"1e", x"1d", x"f0", x"f7", x"f1", x"fe", x"15",
    x"08", x"fa", x"03", x"ff", x"05", x"f9", x"fb", x"04",
    x"01", x"04", x"06", x"00", x"ff", x"fd", x"06", x"04",
    x"00", x"04", x"e5", x"d8", x"e7", x"9f", x"ba", x"e2",
    x"ca", x"9f", x"bb", x"44", x"10", x"19", x"0c", x"00",
    x"f0", x"01", x"cb", x"bc", x"22", x"0a", x"12", x"1c",
    x"11", x"15", x"03", x"06", x"18", x"1d", x"ec", x"04",
    x"fc", x"eb", x"17", x"45", x"37", x"13", x"28", x"50",
    x"49", x"2d", x"23", x"37", x"19", x"fb", x"2f", x"2a",
    x"36", x"27", x"35", x"16", x"05", x"d5", x"f9", x"de",
    x"26", x"18", x"12", x"d7", x"f2", x"c0", x"ca", x"85",
    x"d0", x"20", x"36", x"1a", x"63", x"46", x"11", x"46",
    x"45", x"3a", x"14", x"22", x"0d", x"cb", x"f9", x"11",
    x"a9", x"d5", x"13", x"11", x"f6", x"db", x"2e", x"39",
    x"0a", x"3e", x"5d", x"3c", x"1c", x"5d", x"4f", x"40",
    x"23", x"44", x"3a", x"17", x"20", x"09", x"09", x"28",
    x"3c", x"e4", x"ff", x"71", x"df", x"f9", x"f6", x"4a",
    x"42", x"c8", x"44", x"3c", x"86", x"26", x"48", x"05",
    x"da", x"ec", x"b2", x"b6", x"c5", x"e6", x"e0", x"f7",
    x"ce", x"d8", x"24", x"c5", x"b5", x"0b", x"db", x"d3",
    x"c9", x"e1", x"f7", x"fa", x"f0", x"ed", x"19", x"f9",
    x"f5", x"28", x"12", x"23", x"1e", x"21", x"04", x"07",
    x"b9", x"f6", x"04", x"03", x"2a", x"96", x"d7", x"ee",
    x"77", x"df", x"b6", x"ed", x"f6", x"0a", x"e1", x"1f",
    x"fe", x"fb", x"e6", x"b4", x"cd", x"e9", x"fd", x"12",
    x"e4", x"dc", x"f4", x"3b", x"c8", x"fd", x"ba", x"e9",
    x"0b", x"c4", x"b7", x"e2", x"d9", x"a2", x"a8", x"c8",
    x"ff", x"09", x"e4", x"f9", x"04", x"fb", x"02", x"0c",
    x"c4", x"03", x"10", x"06", x"f5", x"2b", x"ed", x"df",
    x"0e", x"30", x"f8", x"20", x"3d", x"20", x"11", x"18",
    x"3e", x"20", x"f7", x"d5", x"ff", x"12", x"81", x"b0",
    x"39", x"ed", x"aa", x"e7", x"f0", x"2c", x"e4", x"0f",
    x"f0", x"1d", x"ea", x"d7", x"fc", x"cd", x"cb", x"e7",
    x"cb", x"e0", x"1e", x"eb", x"f8", x"f9", x"07", x"3e",
    x"ea", x"07", x"2e", x"d5", x"d7", x"fc", x"dc", x"e8",
    x"fc", x"f3", x"e9", x"02", x"fd", x"0a", x"0e", x"bd",
    x"f2", x"ff", x"f5", x"dc", x"21", x"01", x"bd", x"2a",
    x"df", x"ef", x"18", x"16", x"0e", x"39", x"26", x"10",
    x"ee", x"02", x"fc", x"05", x"05", x"fd", x"02", x"00",
    x"04", x"05", x"ec", x"fb", x"1b", x"22", x"f5", x"fc",
    x"2c", x"27", x"21", x"e6", x"e8", x"0b", x"13", x"01",
    x"1d", x"3b", x"f3", x"df", x"e4", x"1a", x"46", x"11",
    x"fa", x"45", x"35", x"f8", x"24", x"f7", x"e8", x"ff",
    x"5f", x"2c", x"1c", x"21", x"4e", x"28", x"c1", x"fe",
    x"25", x"e8", x"e6", x"13", x"fb", x"10", x"0e", x"3e",
    x"ff", x"02", x"05", x"fc", x"0d", x"e0", x"fc", x"e6",
    x"14", x"ed", x"18", x"dc", x"99", x"df", x"0c", x"d1",
    x"c9", x"ca", x"f3", x"0e", x"2f", x"08", x"e2", x"2b",
    x"00", x"04", x"e2", x"0a", x"f8", x"04", x"0c", x"f9",
    x"52", x"37", x"1b", x"05", x"fd", x"01", x"fe", x"05",
    x"fc", x"fb", x"fe", x"ff", x"d5", x"db", x"fc", x"1d",
    x"fd", x"00", x"12", x"00", x"fb", x"c5", x"d7", x"1e",
    x"d7", x"d9", x"b9", x"e5", x"f8", x"b5", x"f7", x"12",
    x"2e", x"aa", x"f2", x"14", x"80", x"01", x"f5", x"eb",
    x"d4", x"d1", x"27", x"12", x"00", x"0a", x"1c", x"11",
    x"e8", x"d9", x"00", x"04", x"ea", x"da", x"11", x"07",
    x"eb", x"fd", x"f1", x"e1", x"26", x"1f", x"f0", x"fa",
    x"f1", x"00", x"db", x"2a", x"31", x"b3", x"c8", x"19",
    x"f2", x"a1", x"25", x"e7", x"fd", x"fb", x"fd", x"df",
    x"ff", x"f5", x"11", x"fd", x"05", x"00", x"02", x"06",
    x"0c", x"0a", x"0d", x"0c", x"10", x"f0", x"00", x"09",
    x"bc", x"ec", x"0c", x"0f", x"fb", x"0a", x"dd", x"ff",
    x"f5", x"b0", x"e4", x"fc", x"e7", x"e0", x"da", x"dd",
    x"f6", x"0f", x"1c", x"c7", x"09", x"b6", x"df", x"03",
    x"04", x"ff", x"fe", x"fe", x"fe", x"01", x"03", x"04",
    x"00", x"ff", x"37", x"2b", x"08", x"12", x"21", x"f8",
    x"f7", x"fd", x"09", x"21", x"16", x"51", x"3f", x"19",
    x"03", x"3d", x"0f", x"de", x"10", x"15", x"f5", x"db",
    x"07", x"2c", x"fe", x"ec", x"e8", x"29", x"0d", x"05",
    x"19", x"0a", x"e7", x"10", x"23", x"f3", x"05", x"12",
    x"16", x"0b", x"2a", x"e0", x"fa", x"f7", x"01", x"07",
    x"36", x"e4", x"ef", x"e9", x"f7", x"f8", x"08", x"1b",
    x"27", x"14", x"f2", x"0e", x"11", x"0b", x"e5", x"0f",
    x"04", x"02", x"fc", x"01", x"ff", x"05", x"02", x"05",
    x"04", x"04", x"fc", x"fd", x"02", x"00", x"ff", x"05",
    x"fc", x"03", x"f5", x"f1", x"cb", x"e2", x"c3", x"de",
    x"de", x"00", x"bf", x"0a", x"0a", x"f3", x"f7", x"f5",
    x"e4", x"06", x"17", x"02", x"d1", x"f1", x"02", x"d5",
    x"c5", x"e9", x"34", x"d7", x"cb", x"0f", x"e5", x"05",
    x"01", x"ef", x"06", x"21", x"55", x"f9", x"fc", x"fa",
    x"00", x"e4", x"08", x"18", x"1f", x"20", x"12", x"fc",
    x"ed", x"25", x"b1", x"ab", x"f3", x"c3", x"ae", x"c5",
    x"a4", x"ee", x"0e", x"af", x"fa", x"2f", x"be", x"0e",
    x"34", x"03", x"3d", x"29", x"29", x"4d", x"1c", x"fc",
    x"33", x"1c", x"e5", x"0c", x"1c", x"14", x"eb", x"f8",
    x"f5", x"d6", x"f3", x"eb", x"03", x"08", x"dc", x"47",
    x"2f", x"1e", x"34", x"58", x"35", x"1d", x"13", x"5a",
    x"32", x"23", x"12", x"24", x"00", x"f5", x"11", x"18",
    x"07", x"18", x"fd", x"46", x"18", x"05", x"f4", x"e4",
    x"28", x"d3", x"f6", x"33", x"d7", x"e8", x"2c", x"ff",
    x"17", x"26", x"f0", x"db", x"0a", x"00", x"18", x"0e",
    x"3d", x"27", x"f6", x"ba", x"cf", x"d8", x"ff", x"19",
    x"05", x"2e", x"20", x"33", x"e9", x"f3", x"1c", x"b6",
    x"8d", x"ac", x"67", x"6e", x"a3", x"16", x"09", x"0a",
    x"f2", x"f8", x"18", x"ed", x"89", x"c2", x"fe", x"fa",
    x"24", x"07", x"e4", x"d0", x"c0", x"dc", x"f9", x"e0",
    x"05", x"ef", x"2b", x"fe", x"1e", x"15", x"fa", x"3a",
    x"f0", x"a5", x"e0", x"a5", x"d4", x"77", x"11", x"df",
    x"de", x"ef", x"e2", x"01", x"35", x"16", x"fa", x"00",
    x"15", x"23", x"e7", x"e3", x"f0", x"02", x"d4", x"d5",
    x"3b", x"f7", x"1f", x"cf", x"df", x"fb", x"25", x"33",
    x"15", x"1d", x"07", x"1f", x"36", x"24", x"08", x"ca",
    x"d9", x"e5", x"39", x"d9", x"e1", x"2b", x"13", x"0a",
    x"23", x"0c", x"f1", x"14", x"c5", x"d6", x"c5", x"26",
    x"1f", x"d3", x"f9", x"d9", x"1e", x"3f", x"0b", x"fa",
    x"bc", x"c0", x"2d", x"fe", x"08", x"d0", x"f1", x"28",
    x"10", x"0c", x"0e", x"0a", x"17", x"01", x"d7", x"a0",
    x"dd", x"2e", x"e9", x"e3", x"dc", x"09", x"26", x"00",
    x"e4", x"d5", x"f1", x"fd", x"2a", x"03", x"e6", x"40",
    x"13", x"12", x"60", x"d4", x"ea", x"33", x"dc", x"e1",
    x"08", x"fe", x"01", x"04", x"01", x"ff", x"fb", x"03",
    x"05", x"02", x"0f", x"2b", x"cc", x"1e", x"e0", x"b9",
    x"11", x"0d", x"27", x"d5", x"f3", x"49", x"12", x"3d",
    x"37", x"fa", x"1f", x"02", x"1f", x"2a", x"19", x"0f",
    x"39", x"44", x"a2", x"af", x"ac", x"02", x"f8", x"c3",
    x"f9", x"14", x"f4", x"08", x"31", x"23", x"1e", x"43",
    x"53", x"ee", x"30", x"3d", x"e8", x"f6", x"16", x"22",
    x"13", x"2c", x"1c", x"0a", x"00", x"3a", x"08", x"21",
    x"30", x"de", x"b2", x"e3", x"cb", x"1b", x"b5", x"f3",
    x"0d", x"32", x"15", x"13", x"f8", x"29", x"32", x"d2",
    x"04", x"9e", x"f5", x"ff", x"fb", x"1a", x"f0", x"df",
    x"41", x"15", x"d3", x"fd", x"fd", x"03", x"04", x"02",
    x"02", x"ff", x"02", x"01", x"d4", x"f3", x"05", x"22",
    x"1d", x"f6", x"44", x"1c", x"07", x"26", x"15", x"14",
    x"a9", x"e2", x"ba", x"0c", x"e9", x"e1", x"d9", x"cf",
    x"b9", x"44", x"07", x"09", x"86", x"9c", x"9a", x"16",
    x"1d", x"fe", x"f7", x"e9", x"cb", x"f4", x"0e", x"d8",
    x"13", x"11", x"20", x"c6", x"b4", x"da", x"fe", x"d3",
    x"e6", x"13", x"10", x"22", x"48", x"23", x"f6", x"06",
    x"ea", x"ce", x"d7", x"c9", x"dd", x"8b", x"dc", x"19",
    x"80", x"b8", x"17", x"49", x"31", x"de", x"10", x"31",
    x"08", x"21", x"38", x"f7", x"fc", x"fa", x"f3", x"fd",
    x"fc", x"ff", x"f2", x"f4", x"00", x"ef", x"06", x"d7",
    x"3a", x"29", x"36", x"ed", x"fc", x"12", x"e2", x"b6",
    x"d1", x"48", x"04", x"e8", x"09", x"23", x"fc", x"28",
    x"25", x"10", x"08", x"1e", x"d1", x"10", x"05", x"17",
    x"ff", x"fc", x"fa", x"01", x"02", x"04", x"02", x"04",
    x"00", x"b0", x"96", x"8a", x"42", x"20", x"fb", x"d0",
    x"01", x"16", x"4b", x"0e", x"fb", x"d0", x"0b", x"09",
    x"f2", x"31", x"ff", x"6f", x"dd", x"c6", x"48", x"17",
    x"16", x"14", x"d7", x"cb", x"a7", x"c6", x"f5", x"03",
    x"fa", x"2e", x"e0", x"f1", x"08", x"f8", x"c5", x"b0",
    x"16", x"02", x"08", x"3b", x"38", x"1b", x"c5", x"4e",
    x"49", x"13", x"e0", x"ed", x"24", x"21", x"1c", x"e8",
    x"04", x"e8", x"23", x"03", x"10", x"fd", x"22", x"4b",
    x"fa", x"00", x"f7", x"0b", x"ff", x"f9", x"06", x"f9",
    x"fb", x"01", x"00", x"0a", x"07", x"ff", x"00", x"fd",
    x"08", x"04", x"26", x"2f", x"5d", x"ae", x"d9", x"09",
    x"17", x"f7", x"f6", x"2d", x"fd", x"c5", x"ed", x"10",
    x"f1", x"f3", x"1c", x"0f", x"e5", x"de", x"23", x"fe",
    x"16", x"09", x"0f", x"e2", x"9f", x"06", x"1e", x"ff",
    x"d8", x"d8", x"e3", x"e7", x"f5", x"fb", x"64", x"53",
    x"1d", x"55", x"37", x"52", x"1f", x"0a", x"d3", x"cf",
    x"f4", x"ce", x"a6", x"92", x"f6", x"ff", x"e0", x"ce",
    x"1d", x"43", x"00", x"d2", x"06", x"10", x"ca", x"f4",
    x"ca", x"03", x"18", x"07", x"f6", x"d2", x"f8", x"0a",
    x"f9", x"8a", x"12", x"d2", x"cf", x"cf", x"ff", x"0f",
    x"1f", x"fd", x"ec", x"1b", x"f5", x"06", x"27", x"ff",
    x"07", x"98", x"f7", x"17", x"41", x"28", x"0e", x"4c",
    x"11", x"12", x"15", x"10", x"0b", x"e0", x"2e", x"2d",
    x"32", x"fd", x"bd", x"05", x"b5", x"63", x"fb", x"f1",
    x"15", x"dd", x"ad", x"e9", x"1e", x"f5", x"12", x"fa",
    x"ef", x"29", x"b0", x"d9", x"c2", x"e1", x"0e", x"d9",
    x"e9", x"e4", x"1d", x"02", x"e7", x"55", x"e2", x"ae",
    x"ba", x"3b", x"f3", x"b6", x"40", x"03", x"05", x"26",
    x"c9", x"fa", x"0b", x"25", x"47", x"01", x"f1", x"fa",
    x"dc", x"dc", x"df", x"f6", x"04", x"0f", x"c7", x"c7",
    x"cd", x"f8", x"15", x"0e", x"eb", x"ec", x"eb", x"24",
    x"37", x"34", x"09", x"f3", x"e8", x"cc", x"04", x"33",
    x"07", x"1a", x"50", x"e3", x"3e", x"22", x"f7", x"f5",
    x"fe", x"f8", x"db", x"da", x"02", x"cb", x"da", x"f2",
    x"e9", x"1b", x"1a", x"17", x"13", x"28", x"0f", x"e0",
    x"f6", x"e5", x"c3", x"16", x"18", x"b9", x"ff", x"09",
    x"0d", x"1d", x"07", x"10", x"ae", x"94", x"db", x"e4",
    x"ea", x"b6", x"ea", x"ed", x"1d", x"ed", x"dc", x"f9",
    x"0a", x"e0", x"84", x"1f", x"39", x"45", x"cd", x"f7",
    x"e3", x"08", x"73", x"b0", x"fa", x"41", x"2c", x"0a",
    x"20", x"21", x"49", x"2f", x"0a", x"02", x"18", x"31",
    x"00", x"df", x"26", x"eb", x"14", x"1c", x"e9", x"e9",
    x"e5", x"16", x"0b", x"18", x"17", x"23", x"0d", x"25",
    x"1e", x"3a", x"46", x"3b", x"17", x"f1", x"d4", x"36",
    x"e4", x"f4", x"08", x"00", x"f4", x"2d", x"89", x"b7",
    x"15", x"04", x"00", x"05", x"fd", x"01", x"00", x"fd",
    x"fe", x"fb", x"d3", x"ff", x"02", x"28", x"44", x"3f",
    x"16", x"13", x"f0", x"e8", x"d4", x"c1", x"bf", x"c1",
    x"c0", x"95", x"a3", x"c1", x"2a", x"29", x"50", x"12",
    x"f9", x"b1", x"39", x"13", x"fd", x"d7", x"f8", x"e4",
    x"30", x"25", x"c9", x"3e", x"e7", x"b6", x"db", x"f9",
    x"fc", x"1e", x"e2", x"d2", x"c4", x"aa", x"5f", x"e3",
    x"11", x"f9", x"de", x"e0", x"bf", x"f6", x"fd", x"de",
    x"27", x"29", x"01", x"a1", x"f2", x"e1", x"c7", x"d8",
    x"e1", x"13", x"3d", x"08", x"ce", x"00", x"a6", x"f2",
    x"14", x"30", x"cd", x"ce", x"b6", x"32", x"e0", x"97",
    x"8f", x"d4", x"17", x"03", x"08", x"08", x"00", x"04",
    x"03", x"fb", x"f9", x"04", x"e6", x"1a", x"25", x"fd",
    x"17", x"1f", x"32", x"0f", x"14", x"1c", x"ff", x"0c",
    x"0e", x"e8", x"e3", x"99", x"d7", x"fc", x"0d", x"0b",
    x"05", x"25", x"e8", x"c0", x"2f", x"0b", x"c1", x"c4",
    x"07", x"18", x"1c", x"0a", x"32", x"1b", x"28", x"c8",
    x"00", x"17", x"35", x"ee", x"17", x"0e", x"dd", x"f2",
    x"ed", x"07", x"d4", x"c8", x"00", x"c6", x"e0", x"f6",
    x"d6", x"d8", x"0e", x"20", x"33", x"dc", x"f2", x"ec",
    x"3f", x"ff", x"ec", x"1e", x"33", x"11", x"33", x"d4",
    x"c5", x"0f", x"f4", x"ef", x"ff", x"03", x"fb", x"fc",
    x"fb", x"04", x"fc", x"ff", x"fa", x"33", x"23", x"ea",
    x"2a", x"01", x"e3", x"20", x"19", x"1c", x"13", x"22",
    x"1f", x"e4", x"f3", x"f1", x"25", x"29", x"0a", x"f9",
    x"0c", x"0c", x"23", x"09", x"fc", x"c4", x"07", x"0c",
    x"fa", x"05", x"00", x"03", x"00", x"fc", x"fe", x"fd",
    x"fe", x"2d", x"e6", x"06", x"05", x"ed", x"df", x"10",
    x"dc", x"ac", x"0c", x"21", x"fb", x"17", x"f9", x"de",
    x"08", x"d4", x"fd", x"2a", x"04", x"d7", x"15", x"8b",
    x"84", x"ff", x"b0", x"c4", x"48", x"42", x"56", x"38",
    x"06", x"03", x"fe", x"09", x"33", x"e2", x"0d", x"18",
    x"ec", x"bb", x"e8", x"d5", x"e8", x"e4", x"d0", x"05",
    x"3e", x"11", x"0c", x"22", x"1f", x"29", x"31", x"db",
    x"ec", x"d4", x"0f", x"28", x"26", x"23", x"16", x"04",
    x"fc", x"fe", x"00", x"fd", x"fb", x"02", x"01", x"01",
    x"fc", x"00", x"ff", x"04", x"02", x"06", x"06", x"01",
    x"05", x"01", x"d5", x"f7", x"ff", x"c9", x"bb", x"de",
    x"e2", x"da", x"d9", x"c3", x"e6", x"04", x"d6", x"10",
    x"1f", x"eb", x"fc", x"e5", x"d4", x"e0", x"12", x"3b",
    x"38", x"23", x"05", x"2d", x"53", x"e6", x"fd", x"0c",
    x"19", x"33", x"2d", x"c3", x"d7", x"6a", x"de", x"f9",
    x"0f", x"25", x"0b", x"01", x"26", x"1a", x"2e", x"eb",
    x"e3", x"e5", x"21", x"0b", x"18", x"fa", x"11", x"28",
    x"fe", x"f5", x"35", x"f7", x"04", x"13", x"a3", x"15",
    x"14", x"f5", x"d0", x"bd", x"0c", x"03", x"ed", x"fd",
    x"ed", x"ae", x"0b", x"14", x"2d", x"06", x"40", x"2a",
    x"d7", x"b5", x"61", x"28", x"1b", x"46", x"2a", x"46",
    x"54", x"e4", x"69", x"10", x"f5", x"5e", x"f2", x"0f",
    x"d1", x"ab", x"f2", x"cb", x"ac", x"d1", x"d9", x"ff",
    x"3e", x"0b", x"22", x"f4", x"ea", x"9e", x"e1", x"d4",
    x"d9", x"2b", x"15", x"03", x"fc", x"f2", x"cd", x"fa",
    x"11", x"30", x"fe", x"24", x"4d", x"bc", x"ff", x"68",
    x"fd", x"35", x"90", x"1b", x"1c", x"04", x"1e", x"4a",
    x"45", x"33", x"26", x"2e", x"1c", x"27", x"38", x"4c",
    x"57", x"33", x"e5", x"f5", x"26", x"19", x"33", x"08",
    x"1f", x"12", x"16", x"fc", x"dc", x"ea", x"13", x"0b",
    x"ec", x"b1", x"cc", x"b0", x"1e", x"0a", x"1e", x"4d",
    x"36", x"29", x"52", x"3c", x"7a", x"e8", x"ef", x"f4",
    x"ef", x"ec", x"c5", x"f2", x"fe", x"e2", x"c7", x"14",
    x"0a", x"e6", x"d8", x"fe", x"6b", x"9d", x"de", x"cf",
    x"d1", x"8d", x"93", x"c0", x"11", x"dd", x"f2", x"32",
    x"01", x"14", x"f0", x"0e", x"01", x"fe", x"35", x"3c",
    x"37", x"ee", x"ec", x"d0", x"1a", x"f2", x"fc", x"1f",
    x"f8", x"2b", x"12", x"22", x"fa", x"8e", x"d4", x"da",
    x"53", x"5c", x"00", x"04", x"fc", x"1f", x"c7", x"06",
    x"0b", x"e6", x"18", x"f8", x"f0", x"00", x"2d", x"f5",
    x"31", x"2a", x"30", x"34", x"38", x"16", x"1d", x"79",
    x"02", x"13", x"28", x"0f", x"fb", x"2c", x"f8", x"d9",
    x"ff", x"c7", x"ab", x"d8", x"bd", x"af", x"b5", x"0c",
    x"02", x"e5", x"35", x"32", x"2b", x"30", x"58", x"60",
    x"d0", x"f3", x"ec", x"02", x"fc", x"e9", x"17", x"c7",
    x"52", x"ff", x"02", x"fc", x"01", x"fb", x"fb", x"05",
    x"fd", x"05", x"3c", x"20", x"15", x"d0", x"db", x"b1",
    x"f3", x"e8", x"e9", x"f6", x"f9", x"18", x"c2", x"e4",
    x"15", x"b0", x"a9", x"3c", x"01", x"35", x"37", x"10",
    x"2c", x"14", x"00", x"10", x"35", x"d8", x"ba", x"bb",
    x"c1", x"dd", x"ed", x"32", x"15", x"1a", x"f6", x"08",
    x"45", x"e1", x"ed", x"f7", x"d9", x"ef", x"33", x"2c",
    x"1f", x"12", x"3f", x"19", x"f9", x"10", x"33", x"56",
    x"26", x"24", x"16", x"01", x"2f", x"00", x"18", x"13",
    x"f2", x"f0", x"03", x"ee", x"20", x"1f", x"f8", x"73",
    x"48", x"1c", x"0f", x"f5", x"e0", x"d3", x"eb", x"02",
    x"6e", x"fd", x"35", x"fe", x"01", x"fb", x"01", x"07",
    x"ff", x"fd", x"ff", x"fc", x"00", x"ea", x"e2", x"21",
    x"12", x"fd", x"ec", x"f4", x"1c", x"1d", x"0b", x"fe",
    x"d9", x"d5", x"dd", x"05", x"1a", x"11", x"db", x"fd",
    x"16", x"fe", x"f7", x"1e", x"e2", x"e8", x"0d", x"f9",
    x"f8", x"e4", x"f6", x"04", x"f2", x"13", x"0a", x"02",
    x"d7", x"33", x"39", x"e5", x"16", x"03", x"e0", x"cb",
    x"6f", x"d8", x"f7", x"ea", x"06", x"05", x"ff", x"2c",
    x"17", x"31", x"ac", x"46", x"1b", x"b3", x"0e", x"10",
    x"9c", x"e1", x"28", x"f8", x"1f", x"23", x"d8", x"1e",
    x"ff", x"f8", x"3d", x"26", x"03", x"fb", x"fe", x"05",
    x"f8", x"02", x"00", x"f2", x"ff", x"14", x"32", x"25",
    x"1f", x"2f", x"33", x"33", x"0f", x"04", x"27", x"22",
    x"0a", x"f0", x"f5", x"f5", x"54", x"f2", x"de", x"0b",
    x"30", x"11", x"83", x"d0", x"db", x"90", x"b9", x"f1",
    x"01", x"03", x"ff", x"00", x"01", x"fd", x"04", x"04",
    x"04", x"37", x"fc", x"1b", x"17", x"02", x"f0", x"1d",
    x"22", x"13", x"f2", x"26", x"20", x"03", x"1c", x"07",
    x"ef", x"fe", x"10", x"ef", x"f9", x"fb", x"1c", x"ff",
    x"e6", x"28", x"32", x"44", x"48", x"37", x"43", x"15",
    x"39", x"27", x"fc", x"19", x"18", x"e3", x"3b", x"53",
    x"0a", x"15", x"06", x"13", x"09", x"fc", x"33", x"64",
    x"e9", x"d2", x"e2", x"a9", x"ff", x"f7", x"df", x"1b",
    x"0d", x"cd", x"11", x"fa", x"ef", x"05", x"f3", x"df",
    x"fe", x"02", x"fc", x"f7", x"fd", x"fa", x"fe", x"00",
    x"fb", x"ff", x"01", x"00", x"fe", x"00", x"fb", x"fe",
    x"00", x"fb", x"fc", x"03", x"2a", x"df", x"16", x"03",
    x"26", x"1b", x"32", x"ef", x"0a", x"c6", x"dd", x"ec",
    x"e8", x"d8", x"c0", x"65", x"ef", x"00", x"04", x"f7",
    x"0e", x"16", x"d8", x"d5", x"09", x"eb", x"04", x"e4",
    x"1c", x"12", x"ff", x"23", x"3c", x"50", x"66", x"10",
    x"ff", x"d4", x"d6", x"ef", x"bc", x"d6", x"e3", x"f1",
    x"fc", x"36", x"01", x"d6", x"e9", x"f3", x"f0", x"f2",
    x"dd", x"17", x"29", x"8f", x"d3", x"f5", x"fc", x"1c",
    x"01", x"16", x"05", x"00", x"41", x"28", x"2f", x"50",
    x"63", x"63", x"0f", x"f3", x"e0", x"ed", x"12", x"18",
    x"e3", x"33", x"ff", x"06", x"d4", x"cb", x"1e", x"19",
    x"1c", x"38", x"1e", x"14", x"34", x"2e", x"2d", x"1b",
    x"89", x"ce", x"42", x"1f", x"28", x"21", x"16", x"0d",
    x"df", x"eb", x"1b", x"03", x"20", x"30", x"fd", x"15",
    x"16", x"09", x"38", x"27", x"1d", x"38", x"32", x"ef",
    x"dc", x"f9", x"0f", x"fe", x"dc", x"e3", x"f2", x"06",
    x"ed", x"0b", x"57", x"11", x"16", x"f7", x"28", x"16",
    x"e4", x"d7", x"ee", x"cb", x"38", x"e9", x"fb", x"07",
    x"fd", x"bd", x"25", x"1d", x"2a", x"07", x"32", x"1d",
    x"f9", x"de", x"fc", x"d8", x"dc", x"fd", x"1f", x"48",
    x"e9", x"f7", x"04", x"05", x"23", x"3c", x"21", x"40",
    x"5b", x"5a", x"72", x"59", x"1e", x"08", x"ed", x"b9",
    x"28", x"fd", x"c7", x"c5", x"9a", x"ce", x"ee", x"fd",
    x"eb", x"d6", x"de", x"d5", x"4e", x"35", x"db", x"00",
    x"ed", x"0f", x"c0", x"d3", x"ae", x"03", x"f2", x"ae",
    x"10", x"02", x"4c", x"f8", x"e5", x"d7", x"e5", x"f6",
    x"fd", x"21", x"ef", x"04", x"03", x"0e", x"20", x"28",
    x"26", x"29", x"18", x"00", x"15", x"3f", x"28", x"3b",
    x"0e", x"06", x"f2", x"0a", x"08", x"1e", x"12", x"16",
    x"1d", x"b3", x"22", x"1a", x"eb", x"0c", x"01", x"46",
    x"3d", x"1a", x"39", x"2b", x"27", x"03", x"08", x"22",
    x"28", x"1f", x"51", x"11", x"f5", x"03", x"4f", x"05",
    x"e9", x"22", x"fc", x"14", x"01", x"fa", x"f1", x"1f",
    x"49", x"3b", x"1d", x"e4", x"ae", x"15", x"d9", x"01",
    x"ed", x"c1", x"ba", x"f2", x"d3", x"d1", x"1d", x"f3",
    x"f6", x"ff", x"00", x"02", x"01", x"fe", x"02", x"fe",
    x"00", x"02", x"26", x"e9", x"f7", x"fb", x"ed", x"19",
    x"dc", x"b9", x"e0", x"fd", x"08", x"e9", x"ee", x"d2",
    x"9e", x"15", x"fb", x"0d", x"0e", x"19", x"0a", x"0f",
    x"0c", x"0b", x"ed", x"ff", x"07", x"fc", x"f0", x"f6",
    x"98", x"b5", x"d7", x"a5", x"a9", x"8f", x"db", x"c0",
    x"cc", x"d7", x"d9", x"e0", x"fc", x"ec", x"16", x"01",
    x"18", x"13", x"12", x"32", x"2b", x"42", x"16", x"ec",
    x"20", x"02", x"0d", x"08", x"53", x"38", x"2d", x"2c",
    x"fd", x"11", x"15", x"12", x"0e", x"ce", x"f1", x"c5",
    x"de", x"fe", x"1e", x"fa", x"10", x"d3", x"c4", x"c5",
    x"fe", x"90", x"86", x"ff", x"04", x"03", x"01", x"07",
    x"02", x"07", x"02", x"0b", x"2c", x"30", x"7c", x"14",
    x"39", x"40", x"dc", x"f4", x"0a", x"ff", x"f4", x"1f",
    x"ce", x"ee", x"01", x"25", x"1a", x"17", x"03", x"fa",
    x"1b", x"12", x"0d", x"26", x"c2", x"03", x"29", x"2b",
    x"39", x"38", x"fe", x"19", x"de", x"04", x"d1", x"0e",
    x"fb", x"01", x"35", x"df", x"0d", x"27", x"2c", x"1d",
    x"dc", x"d6", x"dc", x"ef", x"09", x"12", x"e8", x"24",
    x"2c", x"37", x"fb", x"dc", x"d0", x"e9", x"dd", x"cd",
    x"af", x"ba", x"f7", x"ec", x"dc", x"f7", x"d8", x"c8",
    x"ea", x"05", x"e6", x"fd", x"00", x"08", x"00", x"fd",
    x"fc", x"fb", x"07", x"05", x"f9", x"c3", x"c6", x"ed",
    x"ce", x"9f", x"a5", x"25", x"ad", x"b4", x"2e", x"56",
    x"52", x"17", x"30", x"32", x"1e", x"ed", x"f7", x"01",
    x"0d", x"3c", x"4d", x"6f", x"5e", x"4c", x"71", x"52",
    x"01", x"01", x"fe", x"fe", x"fd", x"fe", x"ff", x"02",
    x"02", x"0b", x"3d", x"3d", x"ee", x"fc", x"f3", x"bf",
    x"d6", x"ef", x"c9", x"07", x"23", x"f7", x"12", x"37",
    x"e9", x"07", x"00", x"50", x"1c", x"25", x"e1", x"0b",
    x"18", x"14", x"35", x"2c", x"25", x"d0", x"de", x"ef",
    x"d4", x"c4", x"d2", x"ee", x"bb", x"d5", x"00", x"fb",
    x"cb", x"e5", x"b2", x"12", x"ed", x"f7", x"fa", x"b5",
    x"0e", x"14", x"00", x"f2", x"e5", x"e2", x"f6", x"11",
    x"f3", x"13", x"f9", x"fe", x"fc", x"da", x"cc", x"d9",
    x"0d", x"02", x"01", x"00", x"01", x"03", x"04", x"01",
    x"03", x"ff", x"fc", x"fc", x"01", x"07", x"01", x"ff",
    x"fc", x"02", x"07", x"12", x"10", x"3a", x"2c", x"0f",
    x"34", x"30", x"f2", x"0b", x"03", x"60", x"02", x"ff",
    x"20", x"02", x"a8", x"99", x"fd", x"ff", x"3e", x"08",
    x"0c", x"02", x"f5", x"e6", x"c2", x"28", x"4f", x"32",
    x"fb", x"f5", x"c1", x"d9", x"9d", x"bf", x"c8", x"eb",
    x"e9", x"d5", x"07", x"13", x"c5", x"aa", x"bc", x"5b",
    x"fc", x"03", x"36", x"ef", x"e6", x"11", x"09", x"ff",
    x"e8", x"f4", x"19", x"df", x"2a", x"4d", x"ee", x"04",
    x"fc", x"09", x"32", x"1f", x"1b", x"f9", x"08", x"3c",
    x"28", x"3b", x"e3", x"10", x"ea", x"0e", x"ff", x"0a",
    x"12", x"fe", x"e3", x"fe", x"ec", x"f4", x"ec", x"d6",
    x"e1", x"00", x"f8", x"0e", x"ff", x"df", x"fe", x"e4",
    x"0d", x"25", x"10", x"19", x"2d", x"18", x"03", x"da",
    x"fe", x"1d", x"36", x"e5", x"27", x"3f", x"08", x"0b",
    x"ee", x"ee", x"f1", x"ec", x"37", x"ef", x"e1", x"05",
    x"f6", x"f3", x"de", x"fb", x"f8", x"0f", x"24", x"31",
    x"29", x"30", x"4f", x"fb", x"06", x"ee", x"28", x"3c",
    x"2a", x"12", x"fa", x"ee", x"06", x"1d", x"0d", x"ef",
    x"d8", x"c8", x"f5", x"03", x"28", x"e9", x"ba", x"c2",
    x"1c", x"13", x"ad", x"e3", x"c5", x"15", x"ee", x"2b",
    x"19", x"1e", x"01", x"15", x"f3", x"f4", x"09", x"f2",
    x"f3", x"ff", x"fd", x"e2", x"49", x"fc", x"ff", x"3e",
    x"2c", x"11", x"d4", x"1d", x"0f", x"fd", x"02", x"d9",
    x"e7", x"1c", x"04", x"08", x"0e", x"36", x"2c", x"c8",
    x"13", x"2a", x"f5", x"f7", x"0f", x"e4", x"fe", x"1d",
    x"d4", x"dc", x"03", x"de", x"d9", x"ea", x"ad", x"d6",
    x"c3", x"d8", x"05", x"18", x"0a", x"18", x"2f", x"fe",
    x"e7", x"23", x"2e", x"32", x"2d", x"f2", x"10", x"00",
    x"15", x"db", x"ae", x"c2", x"d5", x"e2", x"00", x"ea",
    x"e3", x"2c", x"07", x"a4", x"ec", x"ae", x"c8", x"36",
    x"e8", x"06", x"fb", x"e7", x"a7", x"16", x"f4", x"33",
    x"0e", x"1c", x"17", x"fe", x"de", x"e1", x"f1", x"0c",
    x"00", x"ee", x"d3", x"d1", x"0e", x"fe", x"11", x"f6",
    x"01", x"0f", x"1f", x"44", x"32", x"23", x"23", x"ec",
    x"f7", x"08", x"34", x"fd", x"10", x"be", x"c3", x"ab",
    x"b4", x"01", x"06", x"01", x"01", x"ff", x"05", x"03",
    x"fd", x"ff", x"1d", x"34", x"4f", x"e9", x"d8", x"cf",
    x"f3", x"ee", x"fb", x"f6", x"ef", x"f6", x"f4", x"e4",
    x"10", x"18", x"11", x"f0", x"07", x"e2", x"2d", x"25",
    x"37", x"28", x"2b", x"01", x"ea", x"21", x"10", x"14",
    x"a3", x"bd", x"7e", x"8c", x"5e", x"66", x"22", x"24",
    x"5e", x"e2", x"e7", x"7e", x"a4", x"a1", x"d6", x"da",
    x"0c", x"30", x"e7", x"fc", x"e5", x"d2", x"d0", x"fa",
    x"0d", x"19", x"3a", x"71", x"f7", x"eb", x"86", x"ca",
    x"d9", x"0e", x"2a", x"0d", x"16", x"2f", x"24", x"ec",
    x"0b", x"c3", x"0e", x"0c", x"39", x"89", x"3b", x"41",
    x"c5", x"fa", x"d8", x"02", x"fb", x"ff", x"02", x"fb",
    x"fa", x"02", x"f8", x"fe", x"09", x"13", x"0f", x"cf",
    x"de", x"ee", x"f1", x"13", x"04", x"23", x"21", x"2f",
    x"39", x"39", x"08", x"17", x"4f", x"0f", x"16", x"fa",
    x"f9", x"19", x"18", x"2c", x"0f", x"1a", x"f9", x"c2",
    x"e9", x"d4", x"14", x"12", x"07", x"26", x"fc", x"e6",
    x"10", x"00", x"ee", x"09", x"f7", x"d4", x"f2", x"e5",
    x"af", x"a9", x"f8", x"02", x"1f", x"27", x"16", x"20",
    x"22", x"18", x"ea", x"00", x"04", x"1c", x"17", x"e3",
    x"2d", x"0b", x"e4", x"f1", x"ed", x"ed", x"05", x"15",
    x"0a", x"e9", x"3b", x"1e", x"02", x"09", x"0c", x"04",
    x"fd", x"ff", x"08", x"fc", x"04", x"09", x"18", x"2b",
    x"11", x"0b", x"1c", x"24", x"26", x"c0", x"5d", x"fc",
    x"f0", x"43", x"f2", x"0b", x"48", x"00", x"e5", x"1f",
    x"0b", x"10", x"f8", x"02", x"15", x"12", x"fc", x"19",
    x"06", x"fb", x"02", x"fc", x"ff", x"00", x"fd", x"fe",
    x"fe", x"2a", x"15", x"0f", x"f9", x"1f", x"0f", x"f9",
    x"1a", x"e4", x"fe", x"ee", x"15", x"ea", x"05", x"04",
    x"f4", x"aa", x"91", x"21", x"03", x"fb", x"25", x"18",
    x"17", x"2e", x"f0", x"06", x"d6", x"fc", x"1b", x"e4",
    x"02", x"03", x"d5", x"0f", x"3d", x"23", x"0c", x"ff",
    x"19", x"13", x"08", x"fa", x"ef", x"c3", x"07", x"1f",
    x"53", x"1a", x"2a", x"f9", x"0b", x"0f", x"08", x"1e",
    x"2a", x"f8", x"1c", x"e0", x"dd", x"c6", x"bb", x"da",
    x"f9", x"01", x"02", x"03", x"ff", x"fb", x"02", x"02",
    x"fe", x"fc", x"02", x"fb", x"fd", x"05", x"ff", x"03",
    x"05", x"02", x"0a", x"dc", x"f4", x"ff", x"09", x"09",
    x"f0", x"fd", x"c1", x"28", x"ff", x"df", x"0d", x"dc",
    x"e4", x"e3", x"e5", x"e8", x"ed", x"05", x"5f", x"ec",
    x"e7", x"08", x"f2", x"03", x"16", x"0e", x"f2", x"c3",
    x"c6", x"aa", x"b3", x"b8", x"cd", x"f5", x"0b", x"f1",
    x"04", x"e6", x"e7", x"1f", x"e0", x"e8", x"ca", x"01",
    x"c6", x"ed", x"31", x"14", x"f4", x"21", x"30", x"35",
    x"34", x"1e", x"2f", x"36", x"1f", x"09", x"ec", x"1c",
    x"ec", x"42", x"24", x"ec", x"28", x"11", x"40", x"31",
    x"df", x"2d", x"1d", x"c8", x"c2", x"19", x"31", x"53",
    x"c4", x"44", x"2d", x"dd", x"c6", x"0b", x"dd", x"a1",
    x"aa", x"ba", x"8b", x"6b", x"2d", x"15", x"00", x"21",
    x"12", x"29", x"29", x"12", x"00", x"01", x"17", x"32",
    x"f6", x"12", x"28", x"f3", x"22", x"51", x"fa", x"ee",
    x"f9", x"fc", x"f1", x"e3", x"fe", x"d0", x"c1", x"16",
    x"8d", x"94", x"14", x"e6", x"d0", x"50", x"06", x"2a",
    x"ff", x"02", x"02", x"fd", x"fa", x"04", x"ff", x"03",
    x"fe", x"fc", x"fe", x"f7", x"03", x"fb", x"fe", x"fa",
    x"fc", x"fe", x"04", x"fb", x"02", x"02", x"fc", x"00",
    x"fb", x"03", x"fb", x"f8", x"f8", x"fd", x"f5", x"fc",
    x"f8", x"fb", x"f8", x"f8", x"02", x"00", x"fc", x"fc",
    x"00", x"ff", x"00", x"03", x"00", x"fe", x"01", x"fb",
    x"fd", x"03", x"03", x"ff", x"ff", x"05", x"ff", x"fb",
    x"fd", x"02", x"fe", x"03", x"01", x"00", x"fd", x"fd",
    x"03", x"00", x"fb", x"00", x"04", x"fc", x"ff", x"02",
    x"03", x"fb", x"00", x"fb", x"fd", x"03", x"fe", x"fb",
    x"00", x"fd", x"fd", x"f7", x"fe", x"03", x"05", x"f6",
    x"01", x"fe", x"01", x"00", x"fd", x"ff", x"fd", x"fe",
    x"01", x"fd", x"fd", x"fe", x"ff", x"fc", x"fc", x"fe",
    x"f6", x"fc", x"fb", x"ff", x"fb", x"fa", x"fa", x"fe",
    x"00", x"f6", x"03", x"ff", x"fa", x"04", x"f8", x"00",
    x"fb", x"f6", x"f7", x"f9", x"fc", x"ff", x"02", x"ff",
    x"00", x"ff", x"01", x"ff", x"00", x"01", x"fc", x"03",
    x"ff", x"03", x"03", x"fb", x"01", x"f9", x"ff", x"00",
    x"00", x"01", x"f9", x"04", x"ff", x"01", x"fc", x"fa",
    x"03", x"02", x"04", x"fc", x"01", x"01", x"05", x"fe",
    x"05", x"05", x"01", x"fb", x"00", x"fd", x"00", x"f7",
    x"fe", x"fa", x"fa", x"01", x"fa", x"01", x"fd", x"fb",
    x"02", x"00", x"fb", x"fb", x"01", x"00", x"fb", x"ff",
    x"00", x"00", x"fc", x"03", x"01", x"01", x"02", x"fb",
    x"04", x"fb", x"00", x"fd", x"fa", x"f9", x"fb", x"00",
    x"fd", x"fb", x"fa", x"fc", x"fa", x"fc", x"fb", x"fb",
    x"fe", x"fa", x"01", x"fd", x"fe", x"ff", x"00", x"00",
    x"00", x"ff", x"fe", x"fc", x"fc", x"fe", x"fb", x"ff",
    x"fe", x"ff", x"f8", x"f6", x"01", x"fb", x"fd", x"fa",
    x"ff", x"fc", x"fb", x"01", x"ff", x"fe", x"ff", x"01",
    x"fa", x"fe", x"fd", x"ff", x"fc", x"fe", x"03", x"04",
    x"01", x"fc", x"04", x"05", x"00", x"fe", x"03", x"03",
    x"fb", x"fb", x"fa", x"ff", x"fc", x"02", x"00", x"fb",
    x"ff", x"04", x"fa", x"fe", x"fb", x"03", x"fe", x"04",
    x"04", x"fd", x"fd", x"fb", x"fd", x"03", x"fa", x"00",
    x"02", x"00", x"02", x"00", x"03", x"fd", x"fc", x"02",
    x"ff", x"fb", x"fc", x"f8", x"fa", x"f9", x"fe", x"03",
    x"01", x"02", x"04", x"00", x"fa", x"fa", x"fe", x"fc",
    x"f9", x"ff", x"fa", x"04", x"fc", x"00", x"ff", x"ff",
    x"00", x"fe", x"03", x"01", x"00", x"00", x"01", x"fe",
    x"ff", x"fc", x"fe", x"00", x"fe", x"fb", x"ff", x"fc",
    x"03", x"ff", x"fc", x"fb", x"04", x"ff", x"01", x"fe",
    x"04", x"03", x"fc", x"03", x"ff", x"fe", x"fa", x"01",
    x"01", x"fc", x"fc", x"fa", x"fb", x"fa", x"fd", x"fb",
    x"ff", x"fc", x"fd", x"00", x"01", x"00", x"fd", x"fa",
    x"03", x"01", x"fa", x"ff", x"02", x"03", x"01", x"ff",
    x"00", x"03", x"03", x"01", x"ff", x"04", x"fd", x"fd",
    x"fe", x"fe", x"fd", x"02", x"01", x"fd", x"fe", x"00",
    x"fc", x"fa", x"fb", x"02", x"fd", x"fe", x"02", x"fe",
    x"00", x"fd", x"fd", x"ff", x"ff", x"fa", x"04", x"ff",
    x"fc", x"fc", x"02", x"02", x"ff", x"04", x"ff", x"f8",
    x"fd", x"00", x"00", x"05", x"01", x"05", x"fc", x"fd",
    x"04", x"fe", x"fc", x"fa", x"00", x"fe", x"fb", x"fb",
    x"f9", x"fd", x"03", x"ff", x"fc", x"01", x"01", x"04",
    x"00", x"00", x"04", x"03", x"fd", x"fe", x"ff", x"01",
    x"ff", x"fe", x"fc", x"03", x"03", x"01", x"ff", x"03",
    x"01", x"fe", x"fe", x"fc", x"03", x"00", x"fe", x"fa",
    x"fb", x"fb", x"ff", x"ff", x"fc", x"fb", x"fc", x"fb",
    x"03", x"fd", x"00", x"01", x"ff", x"fc", x"fe", x"04",
    x"fd", x"fa", x"03", x"fd", x"fc", x"fa", x"fe", x"f9",
    x"fe", x"ff", x"fa", x"fe", x"f8", x"00", x"02", x"fe",
    x"fd", x"00", x"fa", x"fb", x"fe", x"f6", x"fe", x"ff",
    x"fc", x"fe", x"01", x"01", x"fd", x"fd", x"fb", x"00",
    x"fb", x"01", x"fe", x"01", x"ff", x"fc", x"f9", x"01",
    x"fd", x"ff", x"fe", x"00", x"00", x"ff", x"fd", x"04",
    x"f7", x"00", x"04", x"fc", x"fb", x"fd", x"01", x"03",
    x"fc", x"03", x"02", x"02", x"01", x"00", x"fc", x"fb",
    x"fc", x"03", x"f8", x"00", x"02", x"ff", x"00", x"03",
    x"fc", x"03", x"ff", x"ff", x"fd", x"fb", x"fb", x"fe",
    x"fd", x"fb", x"ff", x"00", x"fd", x"04", x"fd", x"00",
    x"02", x"01", x"fd", x"fb", x"fe", x"00", x"02", x"01",
    x"fb", x"06", x"fc", x"01", x"02", x"ff", x"fb", x"00",
    x"ea", x"0f", x"06", x"e3", x"f4", x"e5", x"e2", x"ca",
    x"be", x"db", x"08", x"ed", x"24", x"18", x"2b", x"7b",
    x"07", x"02", x"26", x"29", x"31", x"f7", x"15", x"16",
    x"14", x"02", x"f5", x"2f", x"02", x"c6", x"06", x"ec",
    x"f8", x"cd", x"d7", x"0a", x"10", x"17", x"fb", x"1e",
    x"27", x"03", x"10", x"04", x"14", x"fe", x"1d", x"37",
    x"e9", x"f9", x"fe", x"02", x"f0", x"d5", x"f6", x"cf",
    x"e1", x"18", x"e5", x"d4", x"c7", x"c8", x"11", x"b6",
    x"ba", x"40", x"ca", x"91", x"e6", x"fc", x"e0", x"a3",
    x"21", x"1c", x"26", x"f9", x"0d", x"1c", x"fe", x"e6",
    x"16", x"e6", x"02", x"37", x"0f", x"1c", x"1d", x"2a",
    x"1a", x"29", x"e1", x"93", x"d4", x"08", x"c3", x"db",
    x"02", x"cb", x"b5", x"b0", x"b1", x"d5", x"eb", x"bd",
    x"a2", x"e4", x"d4", x"b8", x"bc", x"f5", x"13", x"3f",
    x"2f", x"0b", x"1b", x"f5", x"05", x"1d", x"21", x"13",
    x"1c", x"2e", x"1c", x"f5", x"f9", x"e2", x"20", x"2e",
    x"fd", x"e3", x"c0", x"b4", x"e4", x"07", x"0b", x"3a",
    x"27", x"07", x"3a", x"4d", x"19", x"1c", x"31", x"f1",
    x"08", x"fe", x"29", x"19", x"25", x"54", x"dc", x"be",
    x"13", x"fc", x"04", x"ff", x"ff", x"fd", x"04", x"00",
    x"fd", x"fe", x"02", x"0a", x"45", x"1e", x"cd", x"bb",
    x"1b", x"f6", x"ec", x"e4", x"eb", x"17", x"d6", x"07",
    x"ff", x"f0", x"00", x"0f", x"23", x"09", x"28", x"2a",
    x"4f", x"4d", x"1e", x"1f", x"ff", x"05", x"fe", x"01",
    x"d0", x"bd", x"f3", x"c9", x"a8", x"76", x"e8", x"d4",
    x"f5", x"e8", x"e2", x"06", x"25", x"e1", x"de", x"f9",
    x"15", x"f3", x"11", x"fa", x"dc", x"16", x"10", x"f4",
    x"0e", x"d1", x"ef", x"42", x"2d", x"25", x"89", x"11",
    x"09", x"30", x"33", x"16", x"6a", x"66", x"41", x"5a",
    x"3a", x"19", x"2b", x"fb", x"22", x"b3", x"82", x"d5",
    x"f1", x"95", x"94", x"fd", x"05", x"fd", x"03", x"04",
    x"09", x"fe", x"08", x"04", x"fd", x"eb", x"10", x"0a",
    x"02", x"03", x"07", x"0d", x"20", x"c9", x"ab", x"d1",
    x"f1", x"f3", x"10", x"0b", x"29", x"0e", x"23", x"10",
    x"0d", x"0f", x"26", x"2c", x"13", x"04", x"04", x"c5",
    x"e1", x"ee", x"0c", x"f9", x"e3", x"1c", x"0b", x"05",
    x"38", x"1b", x"03", x"04", x"15", x"d4", x"bf", x"b5",
    x"88", x"ee", x"ed", x"0a", x"0f", x"37", x"14", x"13",
    x"19", x"24", x"f4", x"04", x"e3", x"0b", x"f7", x"e8",
    x"00", x"3f", x"15", x"0a", x"20", x"0b", x"a9", x"f6",
    x"e7", x"f8", x"06", x"f3", x"fe", x"ff", x"07", x"04",
    x"03", x"05", x"05", x"02", x"00", x"cf", x"f3", x"06",
    x"15", x"00", x"f0", x"ff", x"19", x"0c", x"55", x"0a",
    x"fe", x"37", x"21", x"13", x"19", x"cc", x"f8", x"2e",
    x"f3", x"12", x"10", x"e1", x"e5", x"fe", x"b4", x"be",
    x"06", x"fb", x"01", x"00", x"fe", x"02", x"00", x"01",
    x"ff", x"46", x"1d", x"0e", x"4c", x"0c", x"06", x"13",
    x"09", x"11", x"0f", x"d6", x"f3", x"04", x"ef", x"f2",
    x"e5", x"b9", x"c1", x"f0", x"e6", x"f0", x"29", x"05",
    x"3c", x"72", x"32", x"31", x"21", x"26", x"0c", x"bd",
    x"07", x"f4", x"f6", x"f9", x"12", x"e6", x"19", x"d5",
    x"27", x"18", x"1f", x"3e", x"26", x"3f", x"1a", x"fc",
    x"35", x"39", x"12", x"1a", x"00", x"fa", x"f8", x"56",
    x"12", x"38", x"15", x"0b", x"0c", x"13", x"ed", x"a0",
    x"fd", x"03", x"ff", x"fa", x"f9", x"fc", x"fa", x"fd",
    x"03", x"fe", x"fd", x"ff", x"03", x"04", x"fe", x"04",
    x"00", x"fb", x"1d", x"f8", x"0d", x"37", x"44", x"32",
    x"2e", x"56", x"39", x"04", x"dd", x"da", x"f1", x"e0",
    x"e8", x"a8", x"b4", x"c6", x"f6", x"0a", x"3c", x"c3",
    x"df", x"0b", x"ce", x"f9", x"f0", x"e3", x"0f", x"35",
    x"ea", x"d7", x"d3", x"e6", x"dc", x"fc", x"02", x"23",
    x"35", x"00", x"c9", x"c2", x"da", x"cc", x"8e", x"d4",
    x"e8", x"f7", x"06", x"d3", x"de", x"e7", x"c9", x"df",
    x"d7", x"de", x"02", x"d4", x"05", x"da", x"fd", x"f5",
    x"12", x"26", x"41", x"1f", x"38", x"29", x"25", x"e6",
    x"35", x"40", x"16", x"60", x"37", x"52", x"3d", x"21",
    x"35", x"f5", x"3f", x"14", x"01", x"0a", x"04", x"b3",
    x"ef", x"2e", x"d8", x"e3", x"1e", x"2b", x"1c", x"2d",
    x"3c", x"06", x"3a", x"1a", x"f5", x"b9", x"d2", x"1c",
    x"cd", x"0f", x"34", x"52", x"3d", x"6d", x"45", x"3a",
    x"34", x"1b", x"04", x"11", x"0f", x"14", x"f1", x"eb",
    x"83", x"cf", x"df", x"99", x"a7", x"45", x"17", x"0d",
    x"ee", x"ca", x"ca", x"ed", x"e1", x"07", x"12", x"ea",
    x"f2", x"1d", x"fa", x"c6", x"cc", x"d1", x"05", x"f1",
    x"dd", x"04", x"42", x"3e", x"4e", x"1d", x"20", x"42",
    x"12", x"fe", x"28", x"eb", x"06", x"ef", x"fd", x"f9",
    x"ea", x"01", x"11", x"cd", x"d2", x"c9", x"da", x"2e",
    x"0f", x"0b", x"2f", x"2d", x"17", x"12", x"0f", x"f6",
    x"04", x"16", x"5a", x"bd", x"43", x"4b", x"29", x"0b",
    x"0b", x"1f", x"00", x"05", x"fa", x"e2", x"e5", x"fc",
    x"e1", x"3a", x"e4", x"fa", x"ff", x"01", x"df", x"0b",
    x"08", x"e7", x"c7", x"e2", x"fc", x"ee", x"3c", x"20",
    x"2d", x"31", x"02", x"25", x"f5", x"ed", x"1a", x"aa",
    x"a1", x"93", x"42", x"f1", x"03", x"f5", x"d7", x"12",
    x"0e", x"16", x"09", x"28", x"ff", x"28", x"2b", x"e7",
    x"c5", x"05", x"b7", x"9f", x"bb", x"07", x"60", x"a7",
    x"e1", x"0b", x"e5", x"19", x"10", x"15", x"18", x"cc",
    x"27", x"34", x"e0", x"2d", x"07", x"04", x"01", x"ba",
    x"05", x"1a", x"03", x"fa", x"13", x"30", x"31", x"3b",
    x"17", x"19", x"37", x"2f", x"24", x"3d", x"17", x"e6",
    x"cc", x"ec", x"f6", x"fd", x"03", x"f6", x"3c", x"44",
    x"2e", x"03", x"02", x"fd", x"01", x"01", x"05", x"fc",
    x"fd", x"03", x"41", x"f1", x"db", x"4e", x"23", x"24",
    x"24", x"0e", x"1d", x"e3", x"ee", x"fa", x"fd", x"f9",
    x"0b", x"a2", x"77", x"c6", x"33", x"2c", x"2c", x"dd",
    x"c9", x"dd", x"9c", x"c8", x"d8", x"d8", x"d2", x"ee",
    x"fd", x"dd", x"c9", x"91", x"18", x"e4", x"01", x"ee",
    x"f6", x"22", x"1f", x"08", x"f8", x"0c", x"ef", x"0d",
    x"e0", x"e7", x"03", x"f5", x"e2", x"1f", x"13", x"10",
    x"fc", x"8c", x"ca", x"e9", x"f4", x"fb", x"bf", x"ec",
    x"02", x"74", x"3b", x"2f", x"5a", x"52", x"04", x"0e",
    x"02", x"05", x"ef", x"f0", x"da", x"fd", x"e7", x"d9",
    x"24", x"e5", x"06", x"02", x"09", x"0d", x"01", x"0c",
    x"09", x"f9", x"00", x"0f", x"f1", x"00", x"25", x"f3",
    x"f8", x"f8", x"da", x"ec", x"e4", x"05", x"02", x"da",
    x"0a", x"e6", x"d7", x"27", x"ef", x"e7", x"37", x"11",
    x"0d", x"14", x"01", x"06", x"01", x"f3", x"ef", x"ec",
    x"e8", x"02", x"e5", x"e5", x"fc", x"e8", x"dc", x"f7",
    x"e9", x"e2", x"cd", x"d8", x"03", x"26", x"00", x"0c",
    x"17", x"15", x"16", x"05", x"20", x"20", x"07", x"d6",
    x"ae", x"a2", x"19", x"38", x"4d", x"15", x"2b", x"36",
    x"06", x"08", x"25", x"e2", x"de", x"fa", x"03", x"00",
    x"ca", x"e3", x"a3", x"b2", x"ff", x"fc", x"fc", x"00",
    x"fd", x"00", x"fb", x"08", x"03", x"31", x"e0", x"ce",
    x"0d", x"fc", x"e2", x"fc", x"0e", x"ef", x"06", x"c2",
    x"da", x"44", x"1f", x"0f", x"20", x"f1", x"1a", x"06",
    x"c6", x"d5", x"ed", x"10", x"f8", x"13", x"18", x"08",
    x"03", x"fd", x"00", x"fb", x"ff", x"fd", x"fd", x"fe",
    x"fb", x"45", x"e9", x"dc", x"35", x"f4", x"f0", x"f8",
    x"ae", x"a8", x"d2", x"98", x"96", x"ac", x"97", x"a9",
    x"dc", x"b9", x"a0", x"25", x"f0", x"df", x"59", x"da",
    x"ed", x"2d", x"af", x"c3", x"9b", x"27", x"0b", x"11",
    x"3d", x"52", x"34", x"4e", x"4f", x"a4", x"b7", x"b2",
    x"d0", x"e3", x"a8", x"01", x"ea", x"ce", x"44", x"e0",
    x"20", x"33", x"3d", x"4d", x"27", x"1f", x"24", x"64",
    x"74", x"45", x"30", x"3c", x"56", x"29", x"2b", x"5d",
    x"fa", x"fc", x"fd", x"04", x"fe", x"fe", x"01", x"f9",
    x"04", x"02", x"01", x"06", x"fe", x"fd", x"01", x"fe",
    x"00", x"03", x"cf", x"22", x"fc", x"e4", x"1f", x"18",
    x"17", x"13", x"27", x"c5", x"b3", x"d7", x"05", x"0c",
    x"0a", x"03", x"09", x"0c", x"32", x"21", x"1c", x"f7",
    x"12", x"40", x"09", x"e1", x"cf", x"0c", x"f7", x"0c",
    x"05", x"0a", x"06", x"0d", x"cf", x"bd", x"38", x"3c",
    x"2a", x"38", x"08", x"f4", x"0f", x"ff", x"17", x"ef",
    x"b9", x"e1", x"27", x"ed", x"ef", x"07", x"f4", x"ff",
    x"0b", x"ba", x"d6", x"cf", x"dc", x"d9", x"d5", x"ec",
    x"01", x"07", x"14", x"15", x"ef", x"c3", x"de", x"00",
    x"e4", x"d9", x"eb", x"1f", x"1f", x"0e", x"2d", x"2b",
    x"c9", x"dc", x"12", x"37", x"1b", x"38", x"44", x"36",
    x"34", x"1d", x"51", x"4c", x"1c", x"1f", x"07", x"d7",
    x"c3", x"ba", x"e5", x"a3", x"75", x"cd", x"e2", x"0a",
    x"ac", x"c7", x"e8", x"c3", x"c8", x"ea", x"16", x"e9",
    x"27", x"f4", x"e2", x"08", x"fb", x"f9", x"23", x"00",
    x"3c", x"00", x"c7", x"08", x"22", x"b5", x"09", x"41",
    x"d8", x"e2", x"c7", x"f8", x"d4", x"9c", x"dd", x"de",
    x"f9", x"14", x"2c", x"2a", x"f9", x"ec", x"c9", x"ea",
    x"fd", x"ed", x"eb", x"d0", x"cb", x"11", x"09", x"01",
    x"f1", x"f8", x"2c", x"d5", x"dd", x"09", x"cf", x"e4",
    x"e6", x"1c", x"e7", x"d4", x"e1", x"fc", x"11", x"e5",
    x"d0", x"f7", x"10", x"20", x"0c", x"11", x"05", x"ad",
    x"08", x"02", x"29", x"f5", x"19", x"0e", x"50", x"2a",
    x"24", x"2c", x"0d", x"0b", x"f6", x"f9", x"05", x"cc",
    x"aa", x"eb", x"24", x"2b", x"29", x"18", x"35", x"15",
    x"d6", x"ee", x"ba", x"10", x"26", x"3d", x"22", x"30",
    x"2d", x"05", x"13", x"1e", x"07", x"e3", x"c7", x"a0",
    x"83", x"6d", x"23", x"17", x"23", x"20", x"07", x"d5",
    x"0c", x"b3", x"dc", x"f1", x"03", x"21", x"0b", x"f9",
    x"ff", x"cb", x"ed", x"e6", x"eb", x"cc", x"f7", x"ee",
    x"ee", x"22", x"04", x"08", x"07", x"e3", x"0b", x"fa",
    x"ff", x"31", x"33", x"1d", x"f8", x"be", x"f5", x"fa",
    x"fa", x"fd", x"0f", x"09", x"16", x"23", x"39", x"f1",
    x"1e", x"3b", x"21", x"08", x"f1", x"03", x"ef", x"04",
    x"12", x"e7", x"a5", x"04", x"f0", x"ac", x"1a", x"21",
    x"0f", x"04", x"fd", x"fd", x"01", x"fe", x"04", x"04",
    x"fd", x"02", x"ea", x"e7", x"01", x"ed", x"43", x"10",
    x"40", x"23", x"24", x"19", x"0a", x"16", x"f3", x"ef",
    x"05", x"e2", x"00", x"d7", x"e1", x"25", x"26", x"57",
    x"fe", x"e7", x"19", x"e5", x"dc", x"dd", x"0a", x"0b",
    x"1a", x"14", x"20", x"2b", x"5c", x"2d", x"e9", x"b3",
    x"c2", x"27", x"cc", x"b9", x"f7", x"ce", x"e4", x"f1",
    x"2b", x"0a", x"d4", x"15", x"46", x"0f", x"5c", x"2d",
    x"3c", x"c8", x"ee", x"89", x"18", x"17", x"12", x"0f",
    x"03", x"10", x"4b", x"19", x"fa", x"f3", x"eb", x"cb",
    x"d0", x"bc", x"21", x"04", x"01", x"2a", x"16", x"20",
    x"1e", x"02", x"0f", x"01", x"01", x"07", x"fa", x"ff",
    x"fe", x"f6", x"00", x"fd", x"42", x"f0", x"c5", x"1e",
    x"1a", x"0f", x"fd", x"07", x"15", x"04", x"db", x"14",
    x"ea", x"ed", x"46", x"02", x"00", x"1e", x"f3", x"cd",
    x"cf", x"f3", x"c0", x"b5", x"da", x"9d", x"90", x"e9",
    x"08", x"16", x"06", x"1a", x"4c", x"28", x"48", x"68",
    x"cf", x"9a", x"e6", x"0e", x"06", x"1f", x"03", x"19",
    x"2d", x"23", x"1b", x"10", x"01", x"f5", x"df", x"cb",
    x"a6", x"d4", x"47", x"ff", x"02", x"30", x"0c", x"21",
    x"54", x"0b", x"10", x"e8", x"2c", x"16", x"29", x"40",
    x"27", x"07", x"ec", x"da", x"01", x"02", x"fe", x"fe",
    x"fc", x"fa", x"fd", x"00", x"fd", x"1a", x"25", x"61",
    x"ff", x"1f", x"14", x"fc", x"03", x"c7", x"27", x"b5",
    x"ca", x"24", x"ef", x"fa", x"fb", x"06", x"25", x"55",
    x"07", x"03", x"21", x"dd", x"ce", x"ed", x"12", x"19",
    x"01", x"04", x"fc", x"04", x"03", x"00", x"fc", x"fc",
    x"ff", x"d9", x"f4", x"f1", x"e8", x"14", x"22", x"fd",
    x"04", x"f9", x"d0", x"15", x"d7", x"36", x"1a", x"14",
    x"ef", x"04", x"32", x"f2", x"1a", x"2c", x"4c", x"d7",
    x"d5", x"f6", x"9d", x"aa", x"06", x"11", x"ee", x"07",
    x"2f", x"5e", x"1a", x"35", x"41", x"d1", x"16", x"d0",
    x"19", x"0a", x"1c", x"0e", x"0d", x"13", x"2c", x"ef",
    x"8b", x"fc", x"18", x"44", x"eb", x"18", x"2b", x"12",
    x"0f", x"fc", x"2b", x"20", x"f4", x"0a", x"28", x"20",
    x"fe", x"fd", x"01", x"00", x"07", x"09", x"fe", x"00",
    x"ff", x"01", x"fa", x"fe", x"fd", x"f9", x"fd", x"ff",
    x"f7", x"03", x"4b", x"0b", x"e3", x"f4", x"05", x"0e",
    x"02", x"3b", x"4e", x"06", x"dd", x"23", x"10", x"f9",
    x"09", x"0f", x"0b", x"45", x"2a", x"0b", x"fe", x"0b",
    x"f9", x"0c", x"1b", x"02", x"0c", x"e4", x"ec", x"09",
    x"ea", x"3a", x"48", x"2a", x"57", x"1a", x"20", x"df",
    x"2e", x"0d", x"20", x"da", x"09", x"08", x"16", x"36",
    x"22", x"fa", x"70", x"35", x"0f", x"0e", x"04", x"19",
    x"e6", x"f1", x"f3", x"ea", x"c5", x"0a", x"b7", x"c6",
    x"fb", x"e8", x"e5", x"bd", x"e7", x"d5", x"a7", x"f3",
    x"b7", x"da", x"f8", x"f1", x"0c", x"ce", x"1b", x"0d",
    x"f5", x"14", x"19", x"f3", x"18", x"30", x"1a", x"1e",
    x"10", x"db", x"12", x"f7", x"17", x"da", x"64", x"15",
    x"e8", x"01", x"d6", x"b2", x"c1", x"20", x"00", x"e9",
    x"10", x"d4", x"ec", x"ea", x"c9", x"cf", x"d0", x"69",
    x"18", x"f4", x"c4", x"9f", x"d3", x"2a", x"27", x"1d",
    x"17", x"1c", x"35", x"00", x"fa", x"0a", x"fb", x"02",
    x"02", x"ff", x"02", x"fc", x"03", x"fe", x"fb", x"ff",
    x"fd", x"fb", x"02", x"03", x"ff", x"03", x"fe", x"04",
    x"fe", x"fa", x"02", x"fe", x"fb", x"fc", x"fe", x"02",
    x"ff", x"fb", x"01", x"f7", x"00", x"f8", x"f8", x"fb",
    x"fd", x"f7", x"fa", x"fc", x"05", x"03", x"fe", x"fe",
    x"03", x"01", x"fd", x"fa", x"01", x"fd", x"00", x"fd",
    x"fb", x"ff", x"01", x"04", x"fe", x"fb", x"fd", x"00",
    x"02", x"00", x"fe", x"03", x"fb", x"fa", x"fc", x"fb",
    x"fa", x"fb", x"fb", x"fc", x"fd", x"00", x"fc", x"fe",
    x"fb", x"fb", x"00", x"fe", x"fa", x"00", x"02", x"fc",
    x"01", x"ff", x"fd", x"fa", x"fc", x"fc", x"ff", x"00",
    x"fb", x"ff", x"fe", x"fa", x"01", x"fb", x"fc", x"ff",
    x"fc", x"03", x"01", x"fe", x"fb", x"fa", x"03", x"03",
    x"fe", x"00", x"fb", x"fb", x"02", x"fe", x"fc", x"fb",
    x"fa", x"fb", x"04", x"ff", x"fc", x"01", x"fe", x"01",
    x"ff", x"01", x"ff", x"fc", x"fc", x"00", x"ff", x"fb",
    x"fb", x"fc", x"fa", x"fc", x"04", x"fd", x"fc", x"03",
    x"03", x"02", x"03", x"fa", x"fe", x"fa", x"fd", x"f9",
    x"ff", x"fe", x"00", x"02", x"fc", x"03", x"04", x"ff",
    x"fd", x"fc", x"05", x"03", x"ff", x"02", x"fd", x"fe",
    x"ff", x"fb", x"fd", x"05", x"03", x"ff", x"fd", x"03",
    x"fd", x"fb", x"fa", x"fe", x"fe", x"fe", x"02", x"fa",
    x"fc", x"ff", x"fd", x"02", x"00", x"00", x"01", x"02",
    x"01", x"f9", x"00", x"fa", x"fb", x"04", x"ff", x"fc",
    x"00", x"fb", x"f9", x"04", x"fb", x"fd", x"fb", x"03",
    x"fd", x"01", x"fd", x"fb", x"03", x"00", x"ff", x"fb",
    x"fd", x"02", x"00", x"fe", x"00", x"fe", x"01", x"f7",
    x"fd", x"fc", x"00", x"fd", x"fc", x"fa", x"fd", x"fd",
    x"ff", x"00", x"04", x"fb", x"ff", x"fd", x"fc", x"03",
    x"fd", x"fb", x"fc", x"03", x"fb", x"fa", x"fd", x"fb",
    x"00", x"04", x"04", x"04", x"03", x"00", x"04", x"ff",
    x"fe", x"05", x"02", x"fd", x"fe", x"03", x"fd", x"02",
    x"03", x"00", x"02", x"fc", x"fd", x"03", x"02", x"fd",
    x"fc", x"04", x"00", x"fd", x"fc", x"fc", x"04", x"fc",
    x"03", x"fe", x"ff", x"fc", x"02", x"00", x"02", x"01",
    x"00", x"00", x"fd", x"02", x"02", x"05", x"ff", x"ff",
    x"03", x"02", x"fe", x"03", x"03", x"00", x"04", x"ff",
    x"00", x"ff", x"ff", x"02", x"fb", x"00", x"fc", x"02",
    x"fc", x"01", x"fe", x"fc", x"01", x"fa", x"fd", x"fa",
    x"fa", x"03", x"fb", x"03", x"fb", x"fc", x"fd", x"04",
    x"fe", x"ff", x"fa", x"02", x"03", x"01", x"ff", x"05",
    x"fc", x"02", x"01", x"02", x"fc", x"fa", x"04", x"ff",
    x"04", x"03", x"f9", x"fb", x"ff", x"00", x"03", x"fe",
    x"00", x"00", x"fa", x"00", x"03", x"ff", x"02", x"f7",
    x"fa", x"00", x"fd", x"01", x"fc", x"fa", x"fc", x"f7",
    x"05", x"fb", x"01", x"01", x"fd", x"02", x"ff", x"fc",
    x"fe", x"fd", x"02", x"fc", x"00", x"00", x"fd", x"00",
    x"fc", x"fa", x"ff", x"fe", x"fc", x"ff", x"fe", x"fe",
    x"02", x"fd", x"ff", x"03", x"02", x"fd", x"fc", x"fb",
    x"fd", x"fb", x"fd", x"fd", x"ff", x"fd", x"fd", x"00",
    x"ff", x"fa", x"fe", x"02", x"fb", x"00", x"05", x"02",
    x"01", x"04", x"fd", x"00", x"fb", x"fd", x"fc", x"ff",
    x"ff", x"fe", x"fb", x"00", x"fe", x"02", x"ff", x"02",
    x"fc", x"05", x"03", x"ff", x"03", x"00", x"04", x"fe",
    x"03", x"fc", x"05", x"02", x"02", x"04", x"ff", x"fb",
    x"ff", x"04", x"05", x"fc", x"ff", x"04", x"fd", x"ff",
    x"00", x"03", x"00", x"fc", x"fd", x"ff", x"fe", x"00",
    x"fa", x"fc", x"f9", x"03", x"fb", x"fd", x"fe", x"02",
    x"fe", x"00", x"fd", x"fd", x"01", x"00", x"ff", x"fa",
    x"03", x"01", x"00", x"fc", x"03", x"fe", x"fe", x"fb",
    x"03", x"fa", x"fa", x"04", x"00", x"ff", x"02", x"00",
    x"fb", x"01", x"fd", x"02", x"fc", x"fe", x"ff", x"fd",
    x"fc", x"03", x"03", x"01", x"04", x"fb", x"04", x"03",
    x"fd", x"02", x"fe", x"fa", x"00", x"fd", x"03", x"04",
    x"04", x"00", x"fe", x"fc", x"ff", x"fe", x"fc", x"03",
    x"03", x"03", x"04", x"00", x"00", x"04", x"02", x"fc",
    x"03", x"fb", x"00", x"fa", x"fd", x"fe", x"ff", x"02",
    x"04", x"fa", x"ff", x"fe", x"fd", x"fa", x"fc", x"ff",
    x"fe", x"00", x"fc", x"fc", x"fa", x"ff", x"ff", x"02",
    x"fb", x"00", x"fb", x"05", x"04", x"fe", x"01", x"02",
    x"fc", x"ff", x"fc", x"03", x"fb", x"fc", x"00", x"01",
    x"fd", x"02", x"ff", x"fa", x"03", x"fe", x"fa", x"ff",
    x"03", x"e9", x"0e", x"02", x"e7", x"d5", x"f8", x"12",
    x"3f", x"44", x"54", x"3b", x"02", x"14", x"47", x"e9",
    x"28", x"3f", x"40", x"16", x"f8", x"fb", x"fc", x"de",
    x"21", x"07", x"e0", x"cf", x"c8", x"d7", x"f2", x"e2",
    x"14", x"27", x"02", x"e7", x"11", x"2e", x"5a", x"1d",
    x"3e", x"35", x"0c", x"0c", x"2e", x"48", x"4c", x"41",
    x"c9", x"e8", x"e6", x"de", x"e0", x"e1", x"ee", x"db",
    x"b8", x"f2", x"04", x"25", x"11", x"2a", x"37", x"40",
    x"04", x"26", x"0e", x"04", x"05", x"f6", x"09", x"33",
    x"0e", x"25", x"21", x"1b", x"11", x"38", x"f7", x"f2",
    x"13", x"fd", x"14", x"fd", x"dd", x"c8", x"e1", x"dc",
    x"b4", x"9c", x"f9", x"26", x"eb", x"d7", x"05", x"01",
    x"e5", x"27", x"3b", x"bf", x"ce", x"c3", x"fa", x"ed",
    x"02", x"bb", x"f0", x"0e", x"32", x"17", x"ff", x"51",
    x"05", x"03", x"5d", x"1a", x"44", x"17", x"20", x"a0",
    x"df", x"dc", x"1c", x"de", x"dc", x"0d", x"38", x"27",
    x"3a", x"ed", x"12", x"fd", x"ed", x"fc", x"ff", x"c8",
    x"cb", x"ed", x"d7", x"ef", x"12", x"f5", x"eb", x"29",
    x"0b", x"20", x"2c", x"bc", x"f2", x"07", x"a5", x"fb",
    x"3d", x"01", x"00", x"02", x"02", x"04", x"ff", x"04",
    x"01", x"fd", x"2d", x"1a", x"1a", x"df", x"f8", x"d8",
    x"fa", x"04", x"10", x"50", x"5a", x"65", x"21", x"4c",
    x"4c", x"a0", x"e5", x"f3", x"cd", x"15", x"5f", x"f2",
    x"fa", x"26", x"16", x"fc", x"e9", x"16", x"1e", x"05",
    x"3e", x"43", x"1c", x"1b", x"62", x"37", x"2d", x"01",
    x"f7", x"23", x"15", x"f1", x"27", x"14", x"20", x"40",
    x"26", x"3a", x"2b", x"39", x"33", x"4c", x"31", x"42",
    x"24", x"1c", x"22", x"62", x"c8", x"e0", x"19", x"e0",
    x"f2", x"f5", x"e8", x"0c", x"d7", x"cf", x"f3", x"c7",
    x"fd", x"e6", x"41", x"27", x"34", x"37", x"30", x"2f",
    x"a7", x"41", x"78", x"01", x"02", x"0a", x"fe", x"07",
    x"04", x"06", x"01", x"ff", x"07", x"1d", x"f5", x"23",
    x"f8", x"09", x"2f", x"17", x"f2", x"f9", x"03", x"e7",
    x"fb", x"eb", x"fd", x"34", x"ea", x"b6", x"06", x"f6",
    x"f4", x"db", x"d2", x"f0", x"03", x"ed", x"dc", x"19",
    x"0f", x"29", x"16", x"fc", x"17", x"0d", x"11", x"27",
    x"16", x"d2", x"c5", x"11", x"c4", x"b4", x"0a", x"f3",
    x"dc", x"34", x"34", x"27", x"f5", x"f9", x"3c", x"ce",
    x"a2", x"ab", x"ea", x"bf", x"b4", x"f9", x"c9", x"cf",
    x"e6", x"e3", x"d4", x"1c", x"0a", x"08", x"ea", x"19",
    x"2f", x"f3", x"28", x"28", x"01", x"06", x"05", x"03",
    x"06", x"06", x"06", x"fc", x"02", x"1c", x"42", x"60",
    x"e4", x"35", x"3e", x"bd", x"1b", x"11", x"48", x"0f",
    x"ff", x"11", x"e9", x"02", x"10", x"ea", x"e0", x"54",
    x"11", x"f0", x"f6", x"fa", x"ed", x"d2", x"05", x"0b",
    x"fa", x"fc", x"00", x"fd", x"05", x"01", x"fe", x"00",
    x"fd", x"85", x"16", x"1a", x"c2", x"0d", x"18", x"0f",
    x"f8", x"1b", x"68", x"41", x"57", x"36", x"3b", x"24",
    x"f9", x"4b", x"4a", x"e4", x"15", x"38", x"0c", x"ec",
    x"ff", x"49", x"10", x"f7", x"3e", x"3f", x"91", x"16",
    x"44", x"3f", x"d3", x"06", x"20", x"6b", x"56", x"48",
    x"41", x"3a", x"2f", x"26", x"26", x"19", x"7c", x"71",
    x"14", x"f2", x"ec", x"04", x"bf", x"e7", x"e3", x"5a",
    x"35", x"3a", x"17", x"fe", x"d3", x"fc", x"16", x"cb",
    x"03", x"02", x"ff", x"03", x"fd", x"04", x"ff", x"04",
    x"00", x"fe", x"fe", x"04", x"fa", x"04", x"fc", x"04",
    x"04", x"fd", x"36", x"14", x"10", x"6f", x"33", x"0e",
    x"29", x"22", x"05", x"1c", x"e9", x"ee", x"0e", x"09",
    x"f9", x"0f", x"f0", x"ee", x"37", x"23", x"22", x"de",
    x"be", x"0c", x"d6", x"b7", x"cb", x"ef", x"df", x"db",
    x"ec", x"f8", x"dc", x"fd", x"f7", x"21", x"33", x"e8",
    x"bd", x"5f", x"1c", x"fb", x"04", x"03", x"fe", x"39",
    x"f2", x"07", x"27", x"f7", x"0c", x"1b", x"12", x"1f",
    x"e6", x"f3", x"00", x"d5", x"d3", x"01", x"ee", x"e8",
    x"ef", x"11", x"11", x"d4", x"f0", x"fa", x"0a", x"21",
    x"31", x"48", x"ec", x"91", x"d5", x"00", x"eb", x"de",
    x"ec", x"e5", x"02", x"cf", x"f3", x"00", x"dd", x"05",
    x"ef", x"f9", x"f3", x"e1", x"1d", x"bc", x"eb", x"27",
    x"4b", x"25", x"ec", x"f2", x"c0", x"44", x"f5", x"fa",
    x"25", x"fb", x"e2", x"cb", x"fd", x"12", x"ec", x"c6",
    x"e7", x"e1", x"b3", x"f0", x"27", x"ff", x"0a", x"ee",
    x"f6", x"e6", x"f5", x"0c", x"e1", x"15", x"03", x"e1",
    x"e6", x"c9", x"de", x"ba", x"b8", x"34", x"01", x"22",
    x"19", x"b2", x"e5", x"d3", x"9d", x"c3", x"e0", x"00",
    x"fd", x"f5", x"2c", x"2d", x"12", x"03", x"07", x"25",
    x"16", x"05", x"00", x"ee", x"fd", x"06", x"11", x"ef",
    x"f5", x"1c", x"32", x"d4", x"0c", x"1a", x"23", x"52",
    x"53", x"28", x"2f", x"55", x"2d", x"13", x"d8", x"e4",
    x"1a", x"f1", x"d3", x"f8", x"cc", x"c6", x"df", x"f9",
    x"e0", x"01", x"fa", x"db", x"0e", x"32", x"34", x"33",
    x"41", x"02", x"03", x"06", x"fc", x"be", x"ba", x"a1",
    x"16", x"1f", x"ee", x"24", x"04", x"fe", x"06", x"da",
    x"e3", x"14", x"06", x"0d", x"b0", x"fb", x"ff", x"26",
    x"27", x"2d", x"06", x"0a", x"26", x"0c", x"12", x"21",
    x"57", x"0f", x"ff", x"14", x"32", x"04", x"e6", x"fa",
    x"11", x"55", x"30", x"25", x"e3", x"ed", x"be", x"13",
    x"1b", x"09", x"29", x"1e", x"31", x"fa", x"f8", x"01",
    x"03", x"04", x"10", x"2f", x"04", x"ed", x"11", x"3b",
    x"16", x"3c", x"1e", x"fe", x"1b", x"1c", x"23", x"ec",
    x"c0", x"e4", x"fe", x"0c", x"d0", x"36", x"dd", x"b5",
    x"1b", x"d5", x"c1", x"0f", x"b6", x"c0", x"ee", x"01",
    x"e0", x"fe", x"00", x"ff", x"fd", x"ff", x"fc", x"ff",
    x"02", x"fe", x"4c", x"1c", x"e4", x"34", x"10", x"0c",
    x"c0", x"c4", x"c0", x"f1", x"f8", x"0e", x"04", x"04",
    x"f4", x"1e", x"00", x"c1", x"dd", x"ab", x"c8", x"0d",
    x"f0", x"c7", x"20", x"19", x"0f", x"fd", x"1e", x"03",
    x"f4", x"02", x"19", x"f7", x"f2", x"e8", x"0e", x"1b",
    x"bd", x"ed", x"cd", x"d4", x"d7", x"eb", x"f4", x"f2",
    x"e9", x"f4", x"fa", x"29", x"2f", x"07", x"17", x"19",
    x"ea", x"cf", x"fa", x"36", x"df", x"04", x"f2", x"48",
    x"31", x"f7", x"28", x"26", x"f7", x"e7", x"e0", x"03",
    x"0d", x"fb", x"11", x"17", x"04", x"29", x"10", x"fe",
    x"d5", x"bd", x"ac", x"01", x"08", x"03", x"05", x"09",
    x"0f", x"ff", x"0c", x"0b", x"0b", x"48", x"01", x"31",
    x"1d", x"29", x"de", x"1a", x"06", x"2f", x"22", x"cd",
    x"fc", x"fb", x"ef", x"bb", x"16", x"14", x"15", x"13",
    x"39", x"35", x"06", x"fe", x"30", x"0d", x"15", x"66",
    x"52", x"17", x"25", x"15", x"2d", x"f3", x"f5", x"eb",
    x"06", x"05", x"27", x"f8", x"32", x"1c", x"d6", x"09",
    x"dc", x"02", x"f9", x"0e", x"f2", x"1e", x"ee", x"e7",
    x"e8", x"fe", x"18", x"41", x"43", x"c6", x"cb", x"ee",
    x"13", x"dd", x"f2", x"b5", x"ab", x"e1", x"f6", x"f2",
    x"0d", x"ca", x"eb", x"ff", x"fd", x"03", x"01", x"00",
    x"02", x"08", x"04", x"04", x"fb", x"0d", x"04", x"2e",
    x"d6", x"bb", x"e1", x"0b", x"c6", x"af", x"f7", x"5a",
    x"47", x"38", x"11", x"03", x"35", x"57", x"35", x"01",
    x"26", x"3a", x"00", x"30", x"31", x"58", x"65", x"72",
    x"fd", x"05", x"02", x"fb", x"03", x"02", x"fc", x"fd",
    x"06", x"04", x"08", x"10", x"10", x"35", x"53", x"1f",
    x"d4", x"ed", x"d4", x"c0", x"ce", x"d9", x"06", x"21",
    x"c9", x"00", x"19", x"6e", x"47", x"44", x"5b", x"10",
    x"0b", x"2a", x"2b", x"1a", x"0d", x"ee", x"0f", x"00",
    x"f7", x"f8", x"cc", x"b4", x"e2", x"07", x"db", x"f1",
    x"cd", x"e5", x"05", x"ca", x"d9", x"01", x"32", x"14",
    x"9c", x"25", x"da", x"d8", x"0c", x"d0", x"e2", x"2b",
    x"28", x"f9", x"12", x"0a", x"f6", x"01", x"12", x"00",
    x"ff", x"0a", x"0a", x"03", x"00", x"04", x"04", x"08",
    x"fe", x"03", x"02", x"02", x"fe", x"06", x"ff", x"f9",
    x"01", x"fe", x"ff", x"e9", x"ea", x"de", x"f3", x"ef",
    x"45", x"49", x"2a", x"1b", x"32", x"1a", x"15", x"20",
    x"f1", x"03", x"e5", x"e8", x"15", x"28", x"2e", x"d8",
    x"ee", x"1d", x"c7", x"e3", x"cf", x"0c", x"08", x"fe",
    x"13", x"40", x"24", x"ed", x"e7", x"f2", x"d0", x"df",
    x"ed", x"d7", x"e0", x"b0", x"aa", x"90", x"d9", x"0e",
    x"ab", x"a9", x"e2", x"e3", x"01", x"f8", x"e0", x"22",
    x"e8", x"e2", x"0d", x"b4", x"d8", x"38", x"09", x"f3",
    x"e7", x"46", x"35", x"3b", x"da", x"24", x"04", x"ea",
    x"19", x"15", x"fe", x"ac", x"ef", x"f2", x"df", x"e9",
    x"2d", x"f8", x"e1", x"1a", x"07", x"fc", x"ec", x"eb",
    x"e9", x"cf", x"9e", x"c0", x"11", x"9d", x"74", x"a9",
    x"b1", x"be", x"e6", x"ed", x"0e", x"01", x"f5", x"ec",
    x"28", x"fe", x"1a", x"98", x"1d", x"30", x"13", x"d7",
    x"01", x"d2", x"fb", x"fe", x"16", x"e3", x"e0", x"0c",
    x"07", x"f7", x"cc", x"ea", x"d1", x"d2", x"a7", x"20",
    x"f8", x"ca", x"c8", x"c8", x"c5", x"e2", x"f4", x"1a",
    x"3b", x"fc", x"1d", x"1d", x"92", x"da", x"15", x"a2",
    x"ff", x"09", x"97", x"05", x"2b", x"de", x"11", x"29",
    x"29", x"25", x"2d", x"d7", x"e8", x"0e", x"1c", x"df",
    x"ef", x"09", x"01", x"c9", x"0d", x"18", x"2e", x"0f",
    x"35", x"25", x"16", x"42", x"2b", x"f2", x"e5", x"c3",
    x"1d", x"eb", x"e5", x"e4", x"19", x"10", x"ee", x"f1",
    x"ef", x"ea", x"0c", x"db", x"e4", x"36", x"22", x"0f",
    x"35", x"10", x"11", x"fe", x"41", x"0d", x"f5", x"22",
    x"20", x"04", x"fe", x"0c", x"28", x"34", x"21", x"1b",
    x"2e", x"13", x"fd", x"09", x"04", x"15", x"fd", x"f0",
    x"ec", x"f1", x"2a", x"36", x"14", x"81", x"3e", x"40",
    x"39", x"54", x"37", x"c7", x"ca", x"ce", x"e6", x"c0",
    x"e9", x"c9", x"1a", x"10", x"a7", x"c6", x"c5", x"da",
    x"be", x"e5", x"e7", x"1a", x"1f", x"0b", x"1d", x"0a",
    x"0d", x"2f", x"01", x"10", x"16", x"0a", x"bf", x"12",
    x"00", x"e8", x"07", x"ea", x"0c", x"02", x"01", x"b3",
    x"b8", x"c9", x"07", x"dc", x"bd", x"16", x"cc", x"de",
    x"fe", x"eb", x"cb", x"e8", x"f8", x"bb", x"99", x"d2",
    x"e1", x"fe", x"03", x"03", x"fd", x"03", x"ff", x"03",
    x"03", x"04", x"18", x"3e", x"1b", x"16", x"ee", x"c7",
    x"0c", x"dc", x"e7", x"fd", x"31", x"4b", x"f2", x"28",
    x"ff", x"f9", x"e3", x"b7", x"b2", x"00", x"45", x"d5",
    x"e2", x"f6", x"20", x"02", x"23", x"39", x"1e", x"04",
    x"3b", x"1c", x"13", x"fe", x"09", x"fd", x"32", x"f5",
    x"c5", x"0b", x"e1", x"bc", x"15", x"3a", x"14", x"17",
    x"1e", x"07", x"0f", x"45", x"21", x"e5", x"23", x"2c",
    x"d2", x"9c", x"ef", x"e5", x"cb", x"f8", x"f2", x"34",
    x"27", x"bf", x"c3", x"28", x"ea", x"0a", x"fa", x"23",
    x"02", x"f7", x"2a", x"31", x"17", x"31", x"1b", x"1f",
    x"ee", x"15", x"2a", x"05", x"06", x"02", x"11", x"06",
    x"04", x"07", x"0b", x"fc", x"66", x"26", x"0d", x"22",
    x"14", x"e8", x"21", x"fc", x"04", x"31", x"24", x"02",
    x"2d", x"3b", x"dd", x"e4", x"b6", x"a0", x"b7", x"e6",
    x"65", x"16", x"fe", x"f4", x"0e", x"08", x"fc", x"20",
    x"3e", x"30", x"0a", x"0c", x"15", x"de", x"f4", x"d1",
    x"d9", x"fb", x"1c", x"d1", x"e5", x"24", x"c4", x"e8",
    x"1e", x"03", x"14", x"e0", x"16", x"10", x"07", x"e2",
    x"05", x"05", x"eb", x"d7", x"cb", x"cc", x"b1", x"e3",
    x"ad", x"ba", x"01", x"da", x"da", x"35", x"e2", x"3c",
    x"01", x"d7", x"fa", x"e1", x"f8", x"f8", x"fb", x"fd",
    x"fa", x"02", x"f2", x"fc", x"05", x"59", x"48", x"8f",
    x"21", x"1f", x"00", x"2d", x"fa", x"f5", x"23", x"1e",
    x"50", x"b9", x"15", x"18", x"21", x"2a", x"1d", x"ee",
    x"eb", x"f7", x"f2", x"d4", x"d9", x"ef", x"e8", x"f1",
    x"04", x"00", x"fe", x"05", x"01", x"04", x"01", x"02",
    x"fe", x"c4", x"f9", x"3b", x"88", x"f9", x"19", x"19",
    x"e3", x"c2", x"06", x"f5", x"f5", x"e1", x"e0", x"0e",
    x"27", x"11", x"e7", x"38", x"49", x"4b", x"5b", x"30",
    x"29", x"3a", x"11", x"06", x"05", x"0e", x"51", x"1c",
    x"2e", x"44", x"eb", x"0d", x"02", x"dd", x"f2", x"0c",
    x"e7", x"01", x"33", x"10", x"25", x"27", x"63", x"e1",
    x"af", x"0a", x"dd", x"9c", x"fa", x"ac", x"bf", x"23",
    x"4c", x"0a", x"1a", x"39", x"ef", x"fe", x"f7", x"df",
    x"03", x"03", x"08", x"08", x"04", x"05", x"02", x"00",
    x"02", x"06", x"04", x"04", x"fd", x"fc", x"fd", x"fb",
    x"07", x"01", x"14", x"07", x"ce", x"f5", x"eb", x"dd",
    x"f8", x"0f", x"0d", x"47", x"07", x"f3", x"24", x"01",
    x"f9", x"17", x"39", x"3c", x"1d", x"3f", x"16", x"20",
    x"32", x"ff", x"d2", x"e8", x"06", x"fe", x"f2", x"e7",
    x"02", x"05", x"f5", x"00", x"dd", x"ee", x"f2", x"92",
    x"8f", x"22", x"01", x"f0", x"07", x"f4", x"cb", x"e9",
    x"a8", x"c3", x"ed", x"de", x"ef", x"b2", x"f6", x"3f",
    x"d3", x"c2", x"fc", x"ce", x"b5", x"ef", x"f7", x"cc",
    x"03", x"0a", x"1b", x"27", x"ff", x"cc", x"1e", x"df",
    x"ef", x"1e", x"da", x"ad", x"dd", x"25", x"c9", x"e8",
    x"0d", x"f9", x"f5", x"07", x"11", x"04", x"dd", x"1c",
    x"f7", x"a5", x"fc", x"28", x"ee", x"de", x"cb", x"c7",
    x"b8", x"9e", x"cc", x"e4", x"ce", x"34", x"3d", x"15",
    x"21", x"f6", x"e2", x"85", x"cb", x"10", x"bd", x"8e",
    x"79", x"d5", x"a7", x"d4", x"d1", x"0e", x"09", x"e7",
    x"e4", x"da", x"e2", x"e0", x"c3", x"f5", x"fa", x"01",
    x"cf", x"cd", x"cf", x"04", x"f9", x"05", x"2f", x"d9",
    x"f8", x"47", x"3d", x"46", x"19", x"14", x"e9", x"ff",
    x"df", x"bd", x"e7", x"c9", x"e4", x"13", x"0f", x"0a",
    x"fc", x"01", x"21", x"09", x"09", x"1f", x"ed", x"15",
    x"20", x"bc", x"a5", x"db", x"0c", x"08", x"2f", x"f2",
    x"fe", x"23", x"10", x"f6", x"cc", x"3d", x"5b", x"be",
    x"f4", x"0b", x"09", x"15", x"30", x"50", x"bb", x"60",
    x"c9", x"06", x"ef", x"fe", x"1c", x"00", x"ff", x"b8",
    x"fa", x"ce", x"39", x"06", x"fe", x"21", x"2b", x"0e",
    x"e0", x"d8", x"93", x"f0", x"e5", x"ac", x"1c", x"09",
    x"c3", x"22", x"36", x"06", x"14", x"fb", x"f9", x"12",
    x"f4", x"d9", x"13", x"17", x"27", x"fd", x"31", x"28",
    x"27", x"48", x"06", x"97", x"d6", x"e1", x"da", x"17",
    x"24", x"f4", x"db", x"fa", x"11", x"bc", x"90", x"33",
    x"cc", x"ca", x"f3", x"da", x"d0", x"cd", x"e7", x"17",
    x"06", x"f5", x"31", x"0f", x"07", x"20", x"18", x"c2",
    x"c9", x"6e", x"be", x"d9", x"b8", x"14", x"25", x"fd",
    x"cd", x"f9", x"f8", x"f3", x"33", x"fa", x"10", x"3f",
    x"2f", x"04", x"cd", x"2f", x"28", x"eb", x"06", x"01",
    x"dc", x"ff", x"fe", x"02", x"fd", x"fd", x"01", x"00",
    x"fd", x"fc", x"2b", x"ef", x"0f", x"c0", x"ad", x"95",
    x"19", x"21", x"31", x"09", x"fb", x"0f", x"0f", x"18",
    x"f2", x"fc", x"e9", x"e0", x"f9", x"12", x"25", x"ff",
    x"2a", x"4d", x"0a", x"ef", x"12", x"f5", x"2d", x"21",
    x"f3", x"06", x"ff", x"2f", x"28", x"23", x"25", x"0b",
    x"06", x"10", x"24", x"e7", x"0a", x"fc", x"ed", x"01",
    x"2b", x"05", x"0b", x"15", x"13", x"39", x"13", x"10",
    x"a7", x"44", x"a0", x"44", x"cd", x"f2", x"71", x"bf",
    x"d9", x"e2", x"f5", x"12", x"ec", x"29", x"39", x"cd",
    x"cf", x"b6", x"ef", x"ed", x"fa", x"24", x"17", x"f0",
    x"2c", x"0b", x"df", x"04", x"fd", x"04", x"fb", x"fd",
    x"fe", x"fb", x"03", x"02", x"3c", x"37", x"cb", x"fd",
    x"f2", x"fe", x"e8", x"0d", x"2c", x"1e", x"35", x"23",
    x"2a", x"3e", x"18", x"16", x"1a", x"e8", x"c0", x"b5",
    x"cc", x"e2", x"e3", x"d3", x"c2", x"f4", x"e6", x"e4",
    x"f4", x"c3", x"f6", x"07", x"23", x"13", x"02", x"06",
    x"d6", x"e4", x"ec", x"22", x"e7", x"0c", x"08", x"02",
    x"09", x"09", x"22", x"19", x"07", x"e8", x"1f", x"1e",
    x"12", x"f1", x"91", x"b5", x"19", x"da", x"12", x"22",
    x"ee", x"18", x"21", x"10", x"b9", x"d5", x"e9", x"29",
    x"1b", x"6a", x"3c", x"f7", x"01", x"f6", x"03", x"fc",
    x"fe", x"02", x"05", x"0c", x"05", x"2a", x"41", x"5c",
    x"24", x"2e", x"51", x"d4", x"26", x"23", x"e6", x"94",
    x"eb", x"d7", x"0b", x"08", x"af", x"99", x"fd", x"c3",
    x"df", x"de", x"fd", x"de", x"d1", x"ae", x"d7", x"ce",
    x"fa", x"02", x"fc", x"fd", x"fe", x"fe", x"02", x"fe",
    x"01", x"d9", x"7e", x"83", x"ee", x"cf", x"c6", x"d6",
    x"1b", x"36", x"98", x"0e", x"14", x"ee", x"06", x"ee",
    x"36", x"0e", x"eb", x"91", x"f5", x"e2", x"db", x"08",
    x"ed", x"2d", x"bc", x"bb", x"0a", x"eb", x"0f", x"eb",
    x"0d", x"1d", x"1f", x"fd", x"10", x"f7", x"12", x"ac",
    x"1c", x"26", x"df", x"35", x"34", x"f9", x"17", x"98",
    x"4f", x"dd", x"d3", x"f4", x"12", x"24", x"16", x"02",
    x"0c", x"bb", x"eb", x"fd", x"c9", x"25", x"0d", x"0f",
    x"02", x"02", x"02", x"08", x"01", x"02", x"02", x"04",
    x"06", x"03", x"fc", x"fe", x"03", x"01", x"fc", x"03",
    x"fd", x"ff", x"13", x"37", x"1d", x"16", x"30", x"19",
    x"e9", x"cc", x"ce", x"22", x"e4", x"d7", x"d9", x"c0",
    x"0b", x"00", x"fd", x"31", x"1e", x"fa", x"dc", x"d9",
    x"07", x"d7", x"2a", x"17", x"df", x"f8", x"e1", x"de",
    x"d4", x"d1", x"ed", x"e8", x"0b", x"0f", x"d5", x"c6",
    x"d6", x"fd", x"e1", x"de", x"e4", x"04", x"09", x"a9",
    x"3c", x"5a", x"17", x"c4", x"a9", x"24", x"07", x"25",
    x"0a", x"ff", x"08", x"33", x"32", x"1b", x"f7", x"bf",
    x"40", x"56", x"f4", x"fe", x"d9", x"ef", x"e9", x"d4",
    x"e4", x"65", x"d3", x"75", x"9d", x"36", x"0e", x"0b",
    x"01", x"43", x"23", x"14", x"07", x"2c", x"fc", x"fa",
    x"2e", x"07", x"38", x"30", x"04", x"af", x"e2", x"bf",
    x"2c", x"ff", x"45", x"13", x"f4", x"fd", x"ff", x"fd",
    x"19", x"34", x"e2", x"5c", x"05", x"d5", x"2b", x"54",
    x"90", x"06", x"99", x"8d", x"0c", x"eb", x"c8", x"05",
    x"02", x"e0", x"dd", x"e7", x"01", x"03", x"1e", x"ff",
    x"9e", x"c6", x"da", x"b4", x"b9", x"e1", x"d7", x"b9",
    x"d1", x"22", x"e9", x"f0", x"2c", x"ea", x"f5", x"06",
    x"fd", x"2f", x"1d", x"1c", x"16", x"20", x"0d", x"35",
    x"1e", x"0d", x"30", x"0b", x"1b", x"f5", x"0b", x"19",
    x"06", x"91", x"b1", x"c9", x"25", x"09", x"e9", x"3a",
    x"29", x"05", x"05", x"19", x"10", x"0d", x"01", x"b8",
    x"c3", x"04", x"34", x"e9", x"27", x"5e", x"b2", x"9a",
    x"e5", x"ac", x"8c", x"f7", x"f0", x"bc", x"fa", x"db",
    x"d9", x"23", x"e0", x"1d", x"0a", x"f3", x"00", x"20",
    x"ab", x"df", x"ca", x"c3", x"d3", x"c2", x"da", x"ee",
    x"f7", x"ec", x"b6", x"bd", x"13", x"12", x"ed", x"42",
    x"27", x"01", x"52", x"1f", x"24", x"49", x"08", x"13",
    x"2b", x"2e", x"2a", x"34", x"4d", x"2d", x"6a", x"45",
    x"31", x"62", x"47", x"30", x"31", x"c3", x"ca", x"d9",
    x"ee", x"0f", x"07", x"f5", x"19", x"19", x"0f", x"1f",
    x"17", x"2c", x"23", x"01", x"2a", x"38", x"0d", x"19",
    x"eb", x"ee", x"fe", x"0d", x"e8", x"e3", x"09", x"33",
    x"e8", x"0f", x"03", x"00", x"f0", x"0f", x"04", x"f1",
    x"c6", x"c8", x"a5", x"e8", x"c7", x"b8", x"1e", x"18",
    x"0b", x"00", x"01", x"fd", x"01", x"fc", x"05", x"04",
    x"ff", x"04", x"fa", x"35", x"1d", x"d7", x"1e", x"15",
    x"0f", x"09", x"2c", x"06", x"e2", x"ca", x"10", x"f0",
    x"db", x"0d", x"0f", x"de", x"25", x"12", x"05", x"f6",
    x"09", x"2f", x"d7", x"12", x"28", x"fa", x"03", x"13",
    x"fb", x"28", x"22", x"22", x"61", x"21", x"ca", x"e6",
    x"fa", x"e6", x"f4", x"ea", x"0e", x"fd", x"f4", x"3b",
    x"04", x"e8", x"24", x"f1", x"f7", x"0b", x"c0", x"de",
    x"e9", x"12", x"19", x"bc", x"f5", x"1b", x"eb", x"d6",
    x"1a", x"09", x"0d", x"da", x"ef", x"fa", x"01", x"c2",
    x"f6", x"fa", x"ef", x"f2", x"da", x"e7", x"f3", x"d6",
    x"fc", x"18", x"2c", x"fa", x"fe", x"04", x"00", x"03",
    x"06", x"fa", x"01", x"02", x"f7", x"05", x"f2", x"df",
    x"ff", x"10", x"02", x"e3", x"e2", x"05", x"da", x"ea",
    x"2f", x"d4", x"d8", x"24", x"c9", x"d9", x"2d", x"3c",
    x"2b", x"07", x"40", x"33", x"e2", x"54", x"40", x"d0",
    x"c8", x"d8", x"d1", x"e7", x"f3", x"fd", x"f6", x"06",
    x"be", x"d9", x"1c", x"d2", x"c9", x"1f", x"b4", x"d7",
    x"3b", x"f8", x"df", x"d0", x"13", x"fa", x"ca", x"27",
    x"f6", x"ef", x"e1", x"1b", x"2b", x"e1", x"05", x"19",
    x"e4", x"1e", x"36", x"68", x"a8", x"2f", x"b6", x"bf",
    x"04", x"11", x"e0", x"cf", x"fc", x"fa", x"07", x"fc",
    x"f5", x"01", x"02", x"03", x"09", x"24", x"ee", x"22",
    x"2f", x"0c", x"08", x"fb", x"ff", x"17", x"d6", x"15",
    x"fa", x"09", x"e9", x"0a", x"cb", x"d0", x"02", x"bf",
    x"ec", x"2c", x"b8", x"f1", x"02", x"85", x"d3", x"10",
    x"01", x"fb", x"ff", x"01", x"fc", x"05", x"fb", x"fc",
    x"fb", x"52", x"32", x"2c", x"45", x"03", x"03", x"31",
    x"02", x"f4", x"ce", x"0c", x"11", x"de", x"07", x"0f",
    x"2f", x"f3", x"bd", x"6d", x"33", x"39", x"3b", x"1d",
    x"2a", x"11", x"fb", x"06", x"e9", x"0f", x"2b", x"0c",
    x"27", x"31", x"1b", x"16", x"f1", x"c9", x"d2", x"06",
    x"df", x"e6", x"d7", x"02", x"eb", x"e8", x"39", x"06",
    x"e0", x"37", x"21", x"c4", x"1d", x"f8", x"f6", x"1a",
    x"04", x"12", x"06", x"1e", x"f0", x"2d", x"33", x"4a",
    x"fc", x"ff", x"0c", x"03", x"07", x"fe", x"ff", x"01",
    x"01", x"ff", x"04", x"ff", x"ff", x"04", x"04", x"05",
    x"00", x"08", x"f9", x"0d", x"fa", x"cd", x"8a", x"9e",
    x"bf", x"65", x"76", x"da", x"df", x"3d", x"e0", x"07",
    x"fb", x"b0", x"0c", x"42", x"4e", x"14", x"f0", x"3a",
    x"0d", x"f8", x"dc", x"1d", x"14", x"14", x"e7", x"ff",
    x"fd", x"fe", x"14", x"2a", x"5d", x"1e", x"f8", x"1e",
    x"27", x"f1", x"e6", x"f7", x"05", x"f9", x"18", x"d6",
    x"bf", x"d3", x"c3", x"00", x"ff", x"cf", x"ed", x"17",
    x"fc", x"ee", x"22", x"2b", x"16", x"e6", x"b8", x"ba",
    x"26", x"14", x"5f", x"2b", x"23", x"09", x"21", x"2c",
    x"25", x"24", x"ae", x"e3", x"ff", x"c5", x"c3", x"1c",
    x"39", x"b0", x"fb", x"13", x"ea", x"fd", x"56", x"15",
    x"2f", x"23", x"5c", x"68", x"39", x"ff", x"02", x"57",
    x"08", x"04", x"27", x"f1", x"e4", x"53", x"11", x"e5",
    x"37", x"da", x"e0", x"40", x"ea", x"de", x"c4", x"f6",
    x"c9", x"c4", x"1e", x"f1", x"d0", x"1a", x"2f", x"b6",
    x"be", x"bc", x"dd", x"02", x"c9", x"c5", x"0b", x"eb",
    x"d5", x"04", x"5d", x"e2", x"cd", x"c3", x"0b", x"fc",
    x"e6", x"15", x"12", x"00", x"4b", x"c4", x"f4", x"15",
    x"e5", x"de", x"02", x"08", x"1b", x"08", x"04", x"0d",
    x"05", x"f8", x"18", x"f5", x"da", x"e9", x"f5", x"ff",
    x"01", x"96", x"81", x"9d", x"0d", x"02", x"f4", x"ef",
    x"f0", x"0f", x"dd", x"e1", x"ea", x"05", x"fc", x"b6",
    x"f2", x"fe", x"0e", x"22", x"16", x"3b", x"10", x"51",
    x"08", x"2b", x"02", x"ef", x"cb", x"b7", x"e3", x"e7",
    x"df", x"49", x"83", x"d7", x"4a", x"21", x"20", x"4a",
    x"c6", x"aa", x"c4", x"e3", x"d7", x"07", x"f9", x"f6",
    x"4d", x"ee", x"0d", x"e9", x"2a", x"31", x"1d", x"0d",
    x"51", x"4a", x"f3", x"2a", x"f9", x"c4", x"fd", x"0b",
    x"5c", x"ec", x"96", x"eb", x"45", x"25", x"fe", x"1b",
    x"2a", x"bd", x"50", x"0e", x"ff", x"e0", x"c1", x"b9",
    x"eb", x"fa", x"02", x"df", x"0d", x"ff", x"12", x"6f",
    x"0d", x"3e", x"44", x"be", x"e0", x"0f", x"dc", x"d1",
    x"f3", x"a4", x"b5", x"ca", x"d3", x"ec", x"0f", x"11",
    x"d8", x"00", x"b2", x"d9", x"f0", x"fa", x"39", x"23",
    x"e5", x"e8", x"e3", x"ef", x"0e", x"fa", x"fd", x"c6",
    x"e6", x"01", x"06", x"03", x"fa", x"ff", x"fc", x"01",
    x"fc", x"01", x"32", x"29", x"2b", x"f0", x"ef", x"06",
    x"28", x"2f", x"30", x"fc", x"01", x"e1", x"f6", x"fa",
    x"14", x"0d", x"07", x"2d", x"22", x"39", x"1a", x"f4",
    x"f9", x"33", x"40", x"e2", x"2e", x"1b", x"da", x"db",
    x"20", x"fd", x"28", x"4a", x"45", x"43", x"53", x"40",
    x"48", x"f8", x"f3", x"02", x"f6", x"b9", x"d4", x"f8",
    x"f1", x"0e", x"04", x"ed", x"07", x"d7", x"c5", x"df",
    x"11", x"74", x"3f", x"e6", x"ec", x"04", x"51", x"bb",
    x"d4", x"ec", x"ff", x"f5", x"3f", x"f4", x"0c", x"3f",
    x"d8", x"a3", x"eb", x"f9", x"f0", x"02", x"12", x"03",
    x"64", x"5b", x"2f", x"0c", x"04", x"fe", x"0a", x"05",
    x"07", x"fc", x"04", x"fb", x"f2", x"d0", x"00", x"f0",
    x"04", x"f0", x"f3", x"fc", x"f8", x"e6", x"e9", x"0b",
    x"32", x"04", x"dc", x"0f", x"02", x"ff", x"f1", x"2d",
    x"2e", x"e8", x"23", x"21", x"8b", x"fe", x"12", x"94",
    x"71", x"9a", x"de", x"ec", x"fd", x"29", x"20", x"39",
    x"c9", x"ff", x"1e", x"f3", x"fa", x"10", x"02", x"bb",
    x"cc", x"ff", x"dd", x"c7", x"1a", x"f3", x"ad", x"37",
    x"0b", x"f9", x"d1", x"39", x"56", x"03", x"e1", x"24",
    x"31", x"e9", x"13", x"02", x"ab", x"f3", x"d4", x"f6",
    x"19", x"18", x"15", x"15", x"ff", x"0a", x"09", x"f4",
    x"fc", x"0b", x"00", x"08", x"08", x"49", x"15", x"ff",
    x"f4", x"0b", x"1a", x"12", x"39", x"f7", x"32", x"d8",
    x"da", x"0b", x"c5", x"fb", x"f1", x"a0", x"f1", x"fb",
    x"35", x"01", x"35", x"f3", x"03", x"2d", x"ad", x"dd",
    x"ff", x"01", x"fd", x"01", x"02", x"02", x"fd", x"fe",
    x"ff", x"54", x"fd", x"fc", x"f3", x"f0", x"ed", x"cd",
    x"e8", x"ef", x"ea", x"0f", x"17", x"1b", x"0e", x"1e",
    x"43", x"0c", x"16", x"5b", x"09", x"1b", x"15", x"19",
    x"f9", x"f8", x"ce", x"e7", x"d4", x"12", x"13", x"0f",
    x"29", x"1c", x"f6", x"32", x"11", x"f1", x"2a", x"31",
    x"1b", x"07", x"0f", x"e0", x"d7", x"dd", x"12", x"49",
    x"2b", x"fd", x"12", x"b5", x"f7", x"14", x"16", x"03",
    x"eb", x"e9", x"0e", x"f3", x"10", x"e8", x"03", x"27",
    x"fd", x"fe", x"fd", x"fd", x"fe", x"fe", x"fe", x"fe",
    x"f9", x"ff", x"fd", x"00", x"07", x"02", x"fe", x"05",
    x"00", x"02", x"07", x"de", x"d8", x"e1", x"ba", x"8c",
    x"fc", x"bd", x"a5", x"25", x"2e", x"f9", x"1e", x"02",
    x"22", x"fe", x"6c", x"bd", x"09", x"f2", x"0a", x"08",
    x"24", x"0e", x"e5", x"fc", x"04", x"f2", x"d6", x"15",
    x"f2", x"05", x"2b", x"49", x"6e", x"5b", x"23", x"11",
    x"09", x"f1", x"f8", x"e8", x"0a", x"22", x"1f", x"2e",
    x"49", x"2c", x"2a", x"ef", x"03", x"33", x"00", x"f5",
    x"0d", x"34", x"48", x"09", x"0a", x"c0", x"f8", x"e9",
    x"07", x"0d", x"19", x"18", x"4f", x"3d", x"19", x"6b",
    x"4c", x"0f", x"57", x"32", x"45", x"00", x"f5", x"20",
    x"a8", x"2c", x"1b", x"14", x"ff", x"02", x"de", x"19",
    x"18", x"64", x"47", x"47", x"09", x"1e", x"13", x"07",
    x"09", x"06", x"6a", x"46", x"25", x"22", x"29", x"21",
    x"4b", x"07", x"16", x"37", x"38", x"18", x"e3", x"11",
    x"04", x"a9", x"08", x"29", x"da", x"0e", x"1a", x"ee",
    x"24", x"23", x"03", x"15", x"d4", x"36", x"0f", x"f9",
    x"02", x"fa", x"fc", x"fb", x"fb", x"fb", x"01", x"f9",
    x"fb", x"fc", x"fc", x"00", x"05", x"fd", x"fc", x"fe",
    x"ff", x"fa", x"02", x"f9", x"fa", x"01", x"f9", x"01",
    x"fc", x"f9", x"f9", x"f5", x"fb", x"ff", x"f4", x"f5",
    x"fe", x"f6", x"fb", x"ff", x"fc", x"00", x"f9", x"ff",
    x"fb", x"ff", x"00", x"f9", x"fd", x"fc", x"fe", x"ff",
    x"ff", x"ff", x"00", x"fa", x"ff", x"fc", x"ff", x"00",
    x"02", x"03", x"fc", x"00", x"05", x"fe", x"fc", x"fe",
    x"fa", x"fb", x"fc", x"fa", x"fd", x"ff", x"fa", x"01",
    x"01", x"02", x"ff", x"fb", x"fd", x"00", x"03", x"f9",
    x"03", x"fd", x"00", x"fb", x"00", x"f9", x"04", x"fd",
    x"f6", x"00", x"ff", x"fd", x"02", x"fb", x"01", x"ff",
    x"fb", x"04", x"f9", x"01", x"fd", x"f9", x"fd", x"fc",
    x"00", x"fe", x"ff", x"fd", x"03", x"02", x"01", x"fc",
    x"00", x"f9", x"00", x"f6", x"00", x"fa", x"01", x"fb",
    x"01", x"fb", x"f9", x"fc", x"00", x"fe", x"ff", x"00",
    x"fc", x"fe", x"f9", x"fd", x"fc", x"fa", x"ff", x"ff",
    x"fa", x"ff", x"ff", x"00", x"00", x"fa", x"00", x"fc",
    x"ff", x"fd", x"fa", x"ff", x"f8", x"02", x"ff", x"fd",
    x"01", x"03", x"00", x"fc", x"04", x"05", x"fc", x"03",
    x"03", x"ff", x"fb", x"fa", x"00", x"fd", x"ff", x"fc",
    x"03", x"fa", x"f9", x"03", x"00", x"00", x"fb", x"fe",
    x"00", x"f9", x"f8", x"00", x"ff", x"fe", x"02", x"03",
    x"fe", x"fc", x"00", x"f9", x"02", x"03", x"fa", x"f7",
    x"fa", x"fc", x"01", x"fa", x"f9", x"ff", x"fc", x"f6",
    x"fd", x"02", x"fc", x"f8", x"00", x"f9", x"04", x"fb",
    x"fe", x"ff", x"fe", x"00", x"f9", x"02", x"01", x"fe",
    x"fa", x"fe", x"fd", x"05", x"ff", x"fd", x"fb", x"02",
    x"fa", x"ff", x"fe", x"fd", x"fb", x"ff", x"fc", x"ff",
    x"fa", x"01", x"fa", x"f7", x"ff", x"fd", x"fc", x"ff",
    x"f8", x"fe", x"fe", x"fd", x"01", x"fb", x"04", x"00",
    x"ff", x"00", x"fe", x"fd", x"01", x"02", x"fc", x"00",
    x"fe", x"fe", x"02", x"fb", x"fe", x"00", x"fe", x"03",
    x"06", x"00", x"05", x"fe", x"00", x"fd", x"ff", x"01",
    x"fc", x"fd", x"fa", x"00", x"fc", x"00", x"ff", x"fa",
    x"fa", x"05", x"01", x"f9", x"fc", x"fe", x"f9", x"fc",
    x"fe", x"04", x"fe", x"01", x"fb", x"01", x"f9", x"fe",
    x"fe", x"fd", x"f9", x"f9", x"fb", x"f5", x"fb", x"fd",
    x"fd", x"fb", x"f8", x"fa", x"00", x"05", x"ff", x"fa",
    x"00", x"06", x"02", x"f9", x"fb", x"ff", x"00", x"fc",
    x"04", x"03", x"01", x"fb", x"ff", x"fc", x"fd", x"04",
    x"05", x"fd", x"ff", x"ff", x"fc", x"f9", x"fd", x"ff",
    x"ff", x"ff", x"fb", x"fa", x"fe", x"02", x"03", x"02",
    x"fe", x"05", x"f9", x"03", x"ff", x"04", x"ff", x"00",
    x"fc", x"fd", x"fb", x"fb", x"fe", x"04", x"02", x"fd",
    x"03", x"ff", x"04", x"fd", x"00", x"01", x"03", x"fd",
    x"fc", x"00", x"05", x"fc", x"00", x"fb", x"fc", x"00",
    x"fe", x"ff", x"fa", x"fd", x"05", x"fa", x"f9", x"fc",
    x"fe", x"f7", x"f9", x"fb", x"ff", x"fc", x"fb", x"fc",
    x"f6", x"ff", x"ff", x"ff", x"02", x"fd", x"fe", x"fc",
    x"00", x"ff", x"ff", x"f8", x"fa", x"fb", x"f9", x"06",
    x"fc", x"fa", x"fc", x"ff", x"fb", x"ff", x"fe", x"ff",
    x"fe", x"02", x"01", x"fa", x"ff", x"fb", x"ff", x"fd",
    x"00", x"ff", x"01", x"f9", x"f9", x"fd", x"fc", x"00",
    x"01", x"fd", x"05", x"fe", x"01", x"05", x"ff", x"05",
    x"ff", x"01", x"fe", x"01", x"fb", x"ff", x"05", x"ff",
    x"03", x"04", x"02", x"fb", x"02", x"fd", x"fc", x"01",
    x"00", x"fc", x"fe", x"ff", x"fa", x"fc", x"01", x"fa",
    x"01", x"fe", x"fd", x"03", x"00", x"f8", x"f9", x"01",
    x"03", x"fb", x"fa", x"fb", x"fd", x"01", x"fa", x"01",
    x"02", x"fc", x"fd", x"f9", x"00", x"00", x"fb", x"04",
    x"fd", x"fc", x"04", x"01", x"01", x"fa", x"01", x"f9",
    x"01", x"03", x"fd", x"05", x"fb", x"fe", x"03", x"01",
    x"fc", x"fb", x"fa", x"05", x"02", x"fd", x"fb", x"00",
    x"fd", x"fd", x"fa", x"fb", x"05", x"ff", x"f9", x"04",
    x"ff", x"fb", x"fb", x"fe", x"fb", x"fb", x"fb", x"fa",
    x"00", x"ff", x"00", x"fb", x"02", x"f9", x"fe", x"00",
    x"f9", x"fa", x"f9", x"ff", x"fd", x"00", x"ff", x"fb",
    x"fd", x"f9", x"fe", x"ff", x"f9", x"03", x"ff", x"00",
    x"04", x"fe", x"fc", x"01", x"06", x"fe", x"fd", x"fe",
    x"fe", x"ff", x"fd", x"fb", x"fd", x"fe", x"fa", x"02",
    x"fe", x"05", x"00", x"fb", x"f9", x"01", x"fe", x"fb",
    x"ef", x"10", x"1b", x"c4", x"ef", x"2a", x"de", x"f5",
    x"ba", x"f3", x"0c", x"fc", x"00", x"ef", x"b1", x"f2",
    x"e7", x"e7", x"c7", x"9c", x"a9", x"f9", x"f8", x"d5",
    x"f7", x"e4", x"ec", x"0c", x"25", x"1c", x"01", x"0d",
    x"1b", x"1a", x"16", x"3d", x"23", x"fe", x"18", x"11",
    x"cb", x"ef", x"05", x"b1", x"d7", x"ce", x"ef", x"0d",
    x"a2", x"d5", x"c1", x"f6", x"14", x"00", x"27", x"2a",
    x"24", x"e8", x"e7", x"15", x"4b", x"26", x"14", x"99",
    x"bf", x"00", x"ec", x"14", x"10", x"22", x"22", x"08",
    x"d2", x"dd", x"f4", x"f2", x"ff", x"52", x"c7", x"fe",
    x"07", x"bc", x"dd", x"a6", x"e4", x"f0", x"f0", x"fa",
    x"03", x"22", x"2b", x"d3", x"12", x"f2", x"62", x"1b",
    x"ee", x"dd", x"d2", x"45", x"46", x"01", x"1e", x"11",
    x"fe", x"1a", x"2a", x"21", x"37", x"1c", x"f4", x"fa",
    x"f2", x"cd", x"19", x"e6", x"a6", x"e0", x"f0", x"fe",
    x"ff", x"f9", x"ed", x"ec", x"04", x"05", x"0e", x"f0",
    x"be", x"c8", x"f2", x"fc", x"45", x"46", x"42", x"fd",
    x"1d", x"0e", x"fa", x"b9", x"ca", x"3c", x"01", x"e0",
    x"2f", x"02", x"c9", x"b0", x"e7", x"fe", x"d5", x"e5",
    x"1b", x"05", x"04", x"ff", x"00", x"01", x"ff", x"04",
    x"04", x"03", x"a3", x"47", x"60", x"c3", x"dd", x"2f",
    x"ee", x"1e", x"38", x"d5", x"21", x"f5", x"c9", x"fc",
    x"f2", x"e1", x"1b", x"0d", x"22", x"02", x"d5", x"12",
    x"28", x"ca", x"f1", x"17", x"09", x"19", x"0f", x"05",
    x"e6", x"0b", x"30", x"ed", x"9a", x"e8", x"e7", x"e2",
    x"f6", x"cd", x"ba", x"e4", x"c9", x"d3", x"d2", x"0b",
    x"2a", x"28", x"ea", x"00", x"36", x"97", x"6e", x"d6",
    x"42", x"44", x"40", x"f8", x"b6", x"fc", x"ef", x"f8",
    x"f1", x"c9", x"fe", x"04", x"d4", x"dd", x"d3", x"14",
    x"e3", x"b6", x"d1", x"06", x"0b", x"ed", x"fc", x"3d",
    x"e7", x"95", x"03", x"05", x"fc", x"04", x"00", x"04",
    x"fc", x"00", x"fe", x"03", x"1e", x"e3", x"c5", x"17",
    x"32", x"27", x"d8", x"e1", x"fd", x"0f", x"0f", x"13",
    x"fc", x"fd", x"fe", x"f9", x"ba", x"f3", x"c6", x"ed",
    x"f1", x"fd", x"06", x"ef", x"63", x"2b", x"f6", x"2f",
    x"ea", x"f5", x"27", x"00", x"11", x"cb", x"1b", x"53",
    x"fc", x"eb", x"f8", x"20", x"eb", x"df", x"d7", x"cf",
    x"28", x"e0", x"d1", x"05", x"d7", x"f8", x"0a", x"f6",
    x"fb", x"06", x"35", x"13", x"e8", x"37", x"29", x"d3",
    x"38", x"44", x"d6", x"f9", x"0b", x"dc", x"c3", x"d0",
    x"08", x"fe", x"b2", x"e9", x"fc", x"f8", x"f8", x"f9",
    x"02", x"00", x"fa", x"01", x"0a", x"14", x"d0", x"eb",
    x"e9", x"e8", x"db", x"d6", x"e4", x"f1", x"fc", x"c0",
    x"c2", x"de", x"02", x"08", x"1a", x"04", x"1f", x"f5",
    x"e1", x"e9", x"d2", x"0c", x"29", x"01", x"f7", x"3c",
    x"02", x"05", x"ff", x"02", x"fd", x"01", x"fe", x"fd",
    x"00", x"e0", x"db", x"d5", x"9f", x"fe", x"f6", x"46",
    x"23", x"12", x"e9", x"e0", x"f8", x"e7", x"22", x"35",
    x"bf", x"14", x"5b", x"23", x"31", x"25", x"f5", x"09",
    x"15", x"24", x"95", x"c2", x"9f", x"c8", x"e6", x"c8",
    x"1a", x"d2", x"ec", x"0b", x"d9", x"f6", x"00", x"19",
    x"22", x"36", x"11", x"de", x"d5", x"e2", x"bc", x"b9",
    x"af", x"cb", x"ee", x"13", x"d5", x"ce", x"e4", x"5d",
    x"11", x"f7", x"fd", x"c5", x"ea", x"ea", x"03", x"fe",
    x"ff", x"03", x"02", x"fd", x"03", x"00", x"02", x"fb",
    x"00", x"fd", x"ff", x"fb", x"fb", x"02", x"fb", x"fe",
    x"00", x"fc", x"14", x"d4", x"c1", x"29", x"fd", x"fd",
    x"0a", x"2b", x"c8", x"19", x"00", x"27", x"22", x"f7",
    x"23", x"c4", x"dd", x"16", x"f1", x"ef", x"e5", x"ab",
    x"ff", x"f8", x"bc", x"f5", x"0b", x"2c", x"2d", x"fd",
    x"37", x"1d", x"3b", x"09", x"c4", x"15", x"14", x"e5",
    x"14", x"e1", x"a0", x"ce", x"e0", x"fc", x"2d", x"6f",
    x"3c", x"31", x"04", x"ef", x"f2", x"24", x"38", x"24",
    x"06", x"18", x"06", x"fe", x"c8", x"d0", x"a8", x"97",
    x"0b", x"33", x"d3", x"de", x"43", x"08", x"ed", x"ad",
    x"c7", x"da", x"da", x"f9", x"ed", x"f7", x"b3", x"be",
    x"2f", x"0b", x"c2", x"d1", x"12", x"d7", x"1c", x"ed",
    x"fd", x"f0", x"1d", x"cf", x"0f", x"e7", x"d1", x"39",
    x"3d", x"f1", x"15", x"e9", x"df", x"34", x"16", x"e3",
    x"f1", x"14", x"18", x"c2", x"db", x"b7", x"24", x"f0",
    x"ff", x"f2", x"0b", x"ef", x"03", x"fa", x"ed", x"05",
    x"06", x"28", x"44", x"f8", x"07", x"fb", x"02", x"f2",
    x"f8", x"3d", x"56", x"f4", x"f3", x"0b", x"fa", x"1e",
    x"5c", x"db", x"be", x"d2", x"58", x"0c", x"f7", x"17",
    x"1a", x"df", x"01", x"0a", x"34", x"0b", x"f4", x"08",
    x"4e", x"16", x"06", x"fe", x"f0", x"ba", x"e1", x"ed",
    x"d7", x"b2", x"75", x"bc", x"37", x"11", x"02", x"3f",
    x"38", x"18", x"2b", x"19", x"1a", x"d3", x"df", x"f6",
    x"fa", x"da", x"03", x"fa", x"ea", x"f8", x"d7", x"bc",
    x"a0", x"e5", x"c3", x"e5", x"36", x"2e", x"41", x"b7",
    x"e1", x"67", x"e8", x"a9", x"13", x"09", x"f2", x"c0",
    x"2f", x"37", x"4d", x"e9", x"2b", x"27", x"e0", x"03",
    x"2a", x"04", x"f8", x"2e", x"2c", x"0f", x"0c", x"25",
    x"3a", x"46", x"cf", x"d2", x"e9", x"0d", x"e3", x"ed",
    x"34", x"51", x"56", x"cc", x"fc", x"27", x"3f", x"32",
    x"f1", x"29", x"4a", x"50", x"f7", x"3d", x"0b", x"1b",
    x"27", x"f8", x"f3", x"1a", x"00", x"37", x"31", x"26",
    x"18", x"fe", x"27", x"fd", x"27", x"45", x"3a", x"fc",
    x"f5", x"0e", x"d3", x"c9", x"12", x"08", x"f5", x"2e",
    x"3c", x"1d", x"51", x"3c", x"04", x"29", x"5d", x"58",
    x"f4", x"0d", x"23", x"e2", x"f1", x"3a", x"fc", x"e0",
    x"f0", x"fb", x"04", x"03", x"00", x"04", x"00", x"fc",
    x"00", x"ff", x"51", x"2a", x"3e", x"0b", x"e1", x"e6",
    x"e7", x"fd", x"cd", x"d5", x"ea", x"23", x"e7", x"e0",
    x"fe", x"13", x"14", x"f7", x"11", x"ed", x"e2", x"f8",
    x"bd", x"fb", x"ff", x"ff", x"f9", x"f5", x"c7", x"fb",
    x"bc", x"a7", x"d5", x"d4", x"a7", x"b1", x"bd", x"d6",
    x"e6", x"c1", x"ba", x"e4", x"ec", x"fe", x"fd", x"48",
    x"15", x"34", x"2b", x"0f", x"e4", x"14", x"03", x"0c",
    x"22", x"3a", x"2b", x"05", x"3a", x"12", x"09", x"c6",
    x"fb", x"12", x"f2", x"f2", x"07", x"f7", x"00", x"fd",
    x"a9", x"0d", x"ef", x"f5", x"11", x"c7", x"a3", x"ea",
    x"d7", x"a0", x"80", x"05", x"03", x"fd", x"05", x"01",
    x"06", x"03", x"09", x"01", x"38", x"22", x"39", x"2b",
    x"16", x"28", x"f7", x"f3", x"3b", x"cd", x"cf", x"c6",
    x"d3", x"bc", x"af", x"fe", x"1b", x"1a", x"37", x"2c",
    x"28", x"26", x"1a", x"0b", x"e4", x"21", x"1d", x"0f",
    x"f9", x"eb", x"dd", x"ea", x"e6", x"f2", x"f1", x"1f",
    x"4a", x"41", x"50", x"ca", x"ed", x"2f", x"03", x"c7",
    x"c0", x"0b", x"fe", x"12", x"20", x"04", x"0f", x"1f",
    x"30", x"46", x"e4", x"fa", x"f3", x"e7", x"da", x"e2",
    x"cc", x"e5", x"e2", x"36", x"21", x"15", x"b6", x"3e",
    x"22", x"b7", x"4f", x"40", x"fb", x"fb", x"fb", x"f9",
    x"01", x"fd", x"f7", x"f7", x"f7", x"18", x"ce", x"d3",
    x"dc", x"d6", x"f4", x"c9", x"b9", x"cf", x"00", x"50",
    x"3b", x"25", x"f7", x"fb", x"c4", x"e8", x"ea", x"11",
    x"32", x"46", x"ff", x"b0", x"ff", x"a6", x"a7", x"c4",
    x"04", x"ff", x"00", x"02", x"06", x"ff", x"fd", x"02",
    x"02", x"17", x"3b", x"41", x"12", x"07", x"21", x"05",
    x"05", x"fc", x"db", x"f2", x"02", x"ef", x"18", x"1b",
    x"01", x"01", x"13", x"33", x"05", x"f4", x"23", x"3b",
    x"23", x"08", x"6d", x"54", x"0e", x"e5", x"cf", x"07",
    x"06", x"d6", x"af", x"d6", x"c9", x"fb", x"f0", x"1c",
    x"dd", x"df", x"f3", x"ed", x"f6", x"3e", x"0c", x"01",
    x"5c", x"ff", x"bf", x"bd", x"07", x"f9", x"da", x"17",
    x"2e", x"d7", x"13", x"0c", x"d2", x"f4", x"f9", x"13",
    x"07", x"fd", x"04", x"f8", x"fc", x"ff", x"fe", x"06",
    x"ff", x"01", x"fc", x"04", x"05", x"00", x"01", x"fe",
    x"01", x"fd", x"c1", x"d8", x"2e", x"eb", x"f8", x"22",
    x"2e", x"07", x"f8", x"04", x"1a", x"2f", x"8c", x"cd",
    x"0c", x"d7", x"85", x"dc", x"10", x"ff", x"02", x"f3",
    x"20", x"14", x"fd", x"1b", x"2a", x"1d", x"36", x"14",
    x"f5", x"cc", x"c0", x"f1", x"fd", x"cf", x"e4", x"06",
    x"08", x"d4", x"04", x"10", x"16", x"08", x"e7", x"04",
    x"09", x"24", x"c5", x"78", x"c9", x"b1", x"e6", x"cf",
    x"8e", x"a4", x"1c", x"bf", x"ab", x"12", x"91", x"55",
    x"bc", x"05", x"1e", x"1f", x"20", x"24", x"48", x"32",
    x"1e", x"63", x"ed", x"28", x"f4", x"f4", x"0d", x"01",
    x"0e", x"10", x"18", x"1d", x"d7", x"06", x"01", x"f9",
    x"1d", x"0b", x"ed", x"db", x"1b", x"5e", x"3a", x"c8",
    x"17", x"19", x"07", x"22", x"18", x"ee", x"f9", x"0d",
    x"1c", x"1c", x"0e", x"28", x"ff", x"1b", x"43", x"54",
    x"4a", x"e9", x"35", x"2d", x"fb", x"fb", x"1f", x"e5",
    x"e1", x"06", x"92", x"df", x"04", x"f3", x"39", x"06",
    x"c8", x"ae", x"f6", x"e4", x"dc", x"ed", x"1e", x"15",
    x"b1", x"28", x"ef", x"0a", x"24", x"20", x"16", x"4d",
    x"48", x"37", x"34", x"2b", x"43", x"02", x"12", x"17",
    x"e2", x"cf", x"a4", x"0e", x"04", x"d7", x"04", x"e3",
    x"b5", x"07", x"02", x"f0", x"45", x"2a", x"25", x"15",
    x"00", x"24", x"29", x"29", x"55", x"03", x"f1", x"b5",
    x"31", x"b2", x"af", x"f1", x"b6", x"c0", x"01", x"05",
    x"0a", x"2f", x"06", x"07", x"eb", x"e7", x"ea", x"14",
    x"aa", x"22", x"00", x"e4", x"09", x"15", x"1f", x"23",
    x"0e", x"e1", x"10", x"ea", x"f7", x"3b", x"30", x"34",
    x"42", x"0b", x"e5", x"f0", x"0a", x"e8", x"03", x"f6",
    x"f6", x"01", x"db", x"d5", x"dd", x"f3", x"b4", x"c4",
    x"31", x"b7", x"f0", x"1d", x"31", x"19", x"88", x"0a",
    x"fd", x"73", x"f9", x"d0", x"dc", x"e3", x"00", x"05",
    x"20", x"1b", x"06", x"20", x"2c", x"1d", x"11", x"34",
    x"32", x"1d", x"7d", x"14", x"11", x"52", x"cf", x"c0",
    x"d6", x"03", x"03", x"1d", x"05", x"07", x"1f", x"d0",
    x"02", x"2a", x"c9", x"d2", x"20", x"0b", x"d4", x"d6",
    x"ba", x"a2", x"a2", x"e9", x"ac", x"91", x"cf", x"de",
    x"fc", x"03", x"fd", x"04", x"00", x"fd", x"00", x"05",
    x"02", x"01", x"7c", x"7d", x"8f", x"22", x"0f", x"f9",
    x"fa", x"f2", x"fc", x"19", x"09", x"ee", x"28", x"fc",
    x"f3", x"11", x"dd", x"ea", x"2b", x"39", x"0e", x"23",
    x"09", x"20", x"04", x"eb", x"05", x"bd", x"c0", x"e5",
    x"c2", x"c5", x"03", x"e6", x"fa", x"35", x"9d", x"a3",
    x"b4", x"c4", x"b1", x"00", x"e6", x"d2", x"19", x"21",
    x"f8", x"ec", x"15", x"f9", x"0b", x"0c", x"28", x"39",
    x"43", x"d2", x"03", x"d2", x"0b", x"2b", x"00", x"1a",
    x"11", x"0b", x"e4", x"d4", x"33", x"0d", x"c4", x"2f",
    x"f3", x"fe", x"39", x"e5", x"d8", x"0f", x"e8", x"cc",
    x"16", x"03", x"15", x"01", x"04", x"03", x"04", x"08",
    x"09", x"0b", x"0d", x"0f", x"33", x"fe", x"23", x"25",
    x"f9", x"26", x"23", x"fa", x"13", x"17", x"ae", x"b3",
    x"0f", x"d7", x"e3", x"d4", x"00", x"fb", x"17", x"22",
    x"43", x"00", x"08", x"f0", x"ef", x"f3", x"04", x"ed",
    x"02", x"e3", x"f0", x"09", x"f9", x"02", x"fd", x"26",
    x"04", x"fb", x"c4", x"ed", x"f9", x"01", x"f4", x"e2",
    x"f3", x"fd", x"05", x"c0", x"1c", x"17", x"eb", x"23",
    x"ee", x"37", x"41", x"3b", x"48", x"4c", x"55", x"3b",
    x"6a", x"32", x"43", x"e5", x"ab", x"f5", x"fe", x"e8",
    x"f6", x"22", x"2a", x"1e", x"ff", x"fe", x"fe", x"fc",
    x"fe", x"fc", x"fe", x"ff", x"07", x"ee", x"a7", x"88",
    x"fb", x"be", x"9b", x"fd", x"f7", x"ce", x"c1", x"88",
    x"99", x"ce", x"c2", x"eb", x"d0", x"00", x"de", x"27",
    x"26", x"3d", x"14", x"f9", x"04", x"e8", x"f7", x"f2",
    x"fc", x"01", x"05", x"00", x"04", x"02", x"ff", x"07",
    x"04", x"26", x"2f", x"4a", x"27", x"f6", x"fe", x"c7",
    x"ee", x"01", x"cc", x"06", x"27", x"d5", x"f8", x"2b",
    x"9e", x"ef", x"0b", x"f7", x"14", x"18", x"77", x"13",
    x"07", x"1a", x"2f", x"32", x"24", x"bc", x"cf", x"fe",
    x"c1", x"ad", x"16", x"09", x"06", x"84", x"a0", x"d1",
    x"b7", x"d4", x"e7", x"fb", x"e8", x"ff", x"49", x"b6",
    x"0e", x"51", x"f4", x"01", x"0f", x"10", x"27", x"4f",
    x"1f", x"f0", x"62", x"1d", x"49", x"20", x"ff", x"f3",
    x"fc", x"fd", x"00", x"02", x"fb", x"fe", x"f9", x"fd",
    x"06", x"fd", x"fe", x"02", x"ff", x"fe", x"f5", x"fd",
    x"fc", x"fc", x"90", x"e4", x"f8", x"fd", x"29", x"2c",
    x"5b", x"0a", x"29", x"f9", x"bd", x"e2", x"fa", x"d7",
    x"29", x"ed", x"03", x"07", x"1c", x"ce", x"d9", x"39",
    x"f2", x"ca", x"16", x"fd", x"ed", x"14", x"2a", x"3d",
    x"16", x"26", x"3d", x"e1", x"1b", x"52", x"db", x"18",
    x"30", x"dd", x"f3", x"e6", x"c8", x"f4", x"2a", x"6d",
    x"23", x"1f", x"26", x"03", x"11", x"ed", x"01", x"f3",
    x"38", x"f0", x"0a", x"13", x"a2", x"c4", x"ea", x"df",
    x"e4", x"f8", x"19", x"1b", x"45", x"21", x"16", x"45",
    x"fe", x"e9", x"c4", x"f7", x"12", x"e8", x"fd", x"f4",
    x"13", x"c1", x"ac", x"30", x"36", x"24", x"12", x"07",
    x"0d", x"f0", x"0e", x"fc", x"e7", x"0c", x"1e", x"be",
    x"e3", x"e7", x"ed", x"f9", x"05", x"0d", x"0f", x"00",
    x"ec", x"1a", x"3a", x"ee", x"2d", x"53", x"d7", x"27",
    x"23", x"a4", x"e6", x"16", x"14", x"fe", x"ff", x"fa",
    x"0b", x"26", x"24", x"35", x"31", x"fe", x"2e", x"58",
    x"0c", x"01", x"0c", x"08", x"fa", x"0d", x"34", x"3a",
    x"2c", x"06", x"cb", x"d5", x"74", x"ea", x"1d", x"a1",
    x"f8", x"05", x"46", x"36", x"33", x"39", x"36", x"2f",
    x"29", x"42", x"41", x"e4", x"ed", x"b4", x"0c", x"e4",
    x"e9", x"18", x"f5", x"0d", x"1c", x"09", x"e9", x"e9",
    x"e6", x"ce", x"cd", x"b5", x"bf", x"28", x"eb", x"c6",
    x"18", x"11", x"24", x"2e", x"1e", x"10", x"e8", x"17",
    x"28", x"27", x"20", x"34", x"23", x"27", x"12", x"ec",
    x"d9", x"13", x"93", x"7a", x"a4", x"de", x"bb", x"cb",
    x"06", x"ac", x"d9", x"fb", x"a9", x"e0", x"e8", x"ff",
    x"f8", x"35", x"1d", x"ee", x"19", x"1d", x"ea", x"1d",
    x"13", x"c9", x"5d", x"e1", x"db", x"48", x"f8", x"da",
    x"fe", x"26", x"e4", x"f7", x"fa", x"25", x"d9", x"01",
    x"23", x"35", x"51", x"3b", x"1d", x"eb", x"0e", x"1f",
    x"29", x"10", x"d1", x"08", x"14", x"fd", x"0c", x"18",
    x"07", x"18", x"ed", x"ef", x"02", x"f5", x"23", x"0c",
    x"02", x"fd", x"f1", x"00", x"03", x"10", x"16", x"03",
    x"d1", x"db", x"f0", x"f2", x"e3", x"e7", x"cf", x"e6",
    x"fb", x"d3", x"dc", x"f9", x"f9", x"ff", x"e1", x"f0",
    x"d6", x"00", x"00", x"fc", x"03", x"01", x"00", x"03",
    x"00", x"03", x"fa", x"e6", x"fc", x"e5", x"bc", x"e1",
    x"dc", x"f8", x"10", x"23", x"13", x"d8", x"38", x"0d",
    x"cb", x"55", x"29", x"34", x"26", x"ec", x"06", x"d0",
    x"d1", x"ab", x"ca", x"83", x"6b", x"1a", x"2b", x"16",
    x"09", x"fc", x"db", x"c4", x"fc", x"39", x"0a", x"16",
    x"1d", x"f9", x"02", x"f2", x"ce", x"ef", x"e1", x"f7",
    x"d5", x"e0", x"f5", x"d9", x"cb", x"dd", x"f9", x"29",
    x"18", x"1b", x"38", x"f4", x"dd", x"17", x"30", x"2b",
    x"20", x"d1", x"ac", x"a9", x"b9", x"c9", x"be", x"e6",
    x"a8", x"99", x"00", x"0d", x"0c", x"02", x"1b", x"00",
    x"14", x"33", x"42", x"00", x"fe", x"06", x"fb", x"f8",
    x"01", x"fe", x"fd", x"05", x"e8", x"df", x"01", x"a8",
    x"78", x"ac", x"a9", x"72", x"98", x"ed", x"09", x"5d",
    x"0d", x"20", x"20", x"1d", x"fc", x"b7", x"16", x"eb",
    x"f0", x"dc", x"d4", x"dc", x"c7", x"c8", x"e0", x"ce",
    x"89", x"98", x"d2", x"a8", x"a4", x"f0", x"d4", x"c3",
    x"3c", x"26", x"0f", x"27", x"29", x"1f", x"29", x"1c",
    x"2f", x"24", x"fe", x"02", x"ed", x"13", x"9d", x"0b",
    x"5a", x"1d", x"02", x"03", x"f9", x"fe", x"f9", x"fa",
    x"fc", x"1d", x"13", x"1c", x"0f", x"cb", x"fe", x"d4",
    x"ae", x"6e", x"c0", x"a3", x"f7", x"02", x"13", x"fb",
    x"fd", x"08", x"fa", x"f0", x"03", x"04", x"e6", x"da",
    x"dc", x"cd", x"cf", x"bf", x"c5", x"8b", x"43", x"21",
    x"0e", x"41", x"00", x"12", x"29", x"15", x"0a", x"0f",
    x"1a", x"1e", x"f7", x"00", x"0f", x"09", x"1e", x"22",
    x"01", x"fe", x"ff", x"04", x"fd", x"fb", x"ff", x"00",
    x"00", x"ef", x"fb", x"d5", x"10", x"f9", x"f2", x"c7",
    x"ed", x"08", x"bc", x"94", x"de", x"a0", x"cb", x"d6",
    x"b0", x"f6", x"53", x"ed", x"c8", x"c3", x"ec", x"e7",
    x"e6", x"bf", x"35", x"2c", x"de", x"ff", x"09", x"12",
    x"11", x"fc", x"fd", x"1a", x"f9", x"c1", x"d8", x"15",
    x"f3", x"0f", x"25", x"d4", x"f8", x"32", x"d4", x"aa",
    x"26", x"04", x"c2", x"fc", x"fd", x"db", x"c6", x"18",
    x"39", x"36", x"25", x"f6", x"36", x"e5", x"06", x"24",
    x"04", x"05", x"ff", x"01", x"02", x"04", x"01", x"04",
    x"05", x"fd", x"fe", x"fd", x"fc", x"03", x"fc", x"04",
    x"01", x"04", x"33", x"2b", x"dd", x"47", x"2a", x"27",
    x"3e", x"39", x"40", x"3f", x"46", x"59", x"48", x"0c",
    x"05", x"22", x"34", x"e9", x"2f", x"3e", x"42", x"0f",
    x"3f", x"34", x"27", x"0e", x"1b", x"e9", x"ff", x"f7",
    x"e2", x"0b", x"e2", x"cf", x"0f", x"15", x"ff", x"fe",
    x"fe", x"d4", x"07", x"29", x"ec", x"26", x"26", x"02",
    x"03", x"3a", x"60", x"2c", x"f9", x"58", x"17", x"b9",
    x"3c", x"ed", x"2e", x"25", x"de", x"f1", x"01", x"d4",
    x"e7", x"d2", x"e1", x"da", x"d6", x"05", x"01", x"eb",
    x"ff", x"26", x"fa", x"30", x"58", x"34", x"19", x"04",
    x"27", x"ff", x"f9", x"18", x"04", x"01", x"f3", x"e7",
    x"db", x"f9", x"1c", x"e8", x"f6", x"d5", x"cc", x"28",
    x"24", x"1f", x"d0", x"f4", x"2d", x"fd", x"fc", x"13",
    x"23", x"dd", x"98", x"ec", x"db", x"c7", x"f9", x"1a",
    x"33", x"d5", x"fa", x"24", x"b7", x"e5", x"2f", x"d4",
    x"d1", x"d0", x"13", x"11", x"16", x"38", x"10", x"1a",
    x"fa", x"04", x"fe", x"fc", x"00", x"01", x"fa", x"02",
    x"00", x"01", x"01", x"fc", x"ff", x"02", x"f8", x"fd",
    x"fd", x"fc", x"03", x"03", x"fe", x"00", x"fb", x"04",
    x"03", x"02", x"01", x"f9", x"fc", x"fc", x"f9", x"f8",
    x"fc", x"fc", x"fb", x"fa", x"03", x"04", x"fc", x"fb",
    x"fe", x"fd", x"ff", x"fc", x"fc", x"fa", x"00", x"fb",
    x"04", x"fe", x"fb", x"00", x"00", x"01", x"fe", x"01",
    x"01", x"fb", x"fd", x"fc", x"04", x"fd", x"ff", x"fb",
    x"fe", x"00", x"ff", x"fc", x"04", x"03", x"02", x"fc",
    x"fb", x"fa", x"04", x"03", x"fa", x"fa", x"02", x"f9",
    x"02", x"00", x"fb", x"ff", x"00", x"fd", x"00", x"fd",
    x"fd", x"f9", x"02", x"03", x"03", x"fd", x"fc", x"fb",
    x"fd", x"fa", x"fb", x"fa", x"fb", x"ff", x"00", x"04",
    x"04", x"fc", x"01", x"00", x"fd", x"fe", x"02", x"02",
    x"fe", x"01", x"fe", x"fc", x"fa", x"f9", x"02", x"02",
    x"f9", x"fd", x"fd", x"02", x"f7", x"fe", x"03", x"02",
    x"04", x"fe", x"fe", x"01", x"fe", x"f9", x"01", x"fd",
    x"fa", x"02", x"00", x"fc", x"fb", x"fa", x"04", x"03",
    x"fe", x"ff", x"01", x"fe", x"fe", x"01", x"fc", x"fc",
    x"fd", x"fd", x"fa", x"fb", x"fd", x"00", x"01", x"02",
    x"05", x"fd", x"02", x"03", x"fc", x"fb", x"fd", x"ff",
    x"fb", x"02", x"fc", x"fc", x"02", x"02", x"fe", x"f7",
    x"01", x"02", x"01", x"ff", x"fd", x"fd", x"fb", x"fe",
    x"04", x"03", x"fe", x"02", x"fa", x"00", x"ff", x"00",
    x"00", x"fb", x"fb", x"fc", x"fd", x"00", x"ff", x"03",
    x"03", x"fc", x"fa", x"01", x"03", x"fb", x"fd", x"00",
    x"fb", x"00", x"f6", x"01", x"03", x"fb", x"fd", x"fe",
    x"fe", x"fb", x"00", x"00", x"fe", x"fa", x"fd", x"03",
    x"fd", x"fb", x"04", x"00", x"fa", x"fd", x"fa", x"fb",
    x"00", x"ff", x"fb", x"fb", x"02", x"fe", x"fb", x"01",
    x"fe", x"ff", x"00", x"03", x"02", x"01", x"04", x"ff",
    x"fe", x"03", x"05", x"05", x"01", x"fe", x"ff", x"f9",
    x"ff", x"fc", x"ff", x"ff", x"fe", x"01", x"01", x"02",
    x"fb", x"04", x"00", x"fd", x"fb", x"fc", x"ff", x"fb",
    x"fc", x"03", x"ff", x"fe", x"00", x"f9", x"00", x"01",
    x"00", x"02", x"00", x"03", x"03", x"01", x"02", x"01",
    x"ff", x"03", x"ff", x"fa", x"04", x"01", x"fe", x"fa",
    x"fe", x"00", x"fe", x"02", x"00", x"02", x"fa", x"fb",
    x"fc", x"fc", x"fe", x"fe", x"01", x"02", x"01", x"fa",
    x"fe", x"03", x"fc", x"fc", x"fd", x"f9", x"fa", x"fc",
    x"01", x"04", x"fb", x"ff", x"03", x"04", x"01", x"04",
    x"00", x"fb", x"00", x"fe", x"fe", x"fc", x"fb", x"fb",
    x"ff", x"ff", x"fb", x"ff", x"fc", x"00", x"fd", x"01",
    x"03", x"01", x"03", x"fc", x"fc", x"fc", x"fe", x"ff",
    x"ff", x"fd", x"f8", x"03", x"fb", x"fc", x"fd", x"f9",
    x"fe", x"ff", x"fd", x"03", x"04", x"fd", x"ff", x"fd",
    x"ff", x"01", x"00", x"fa", x"fd", x"fb", x"02", x"fa",
    x"f7", x"f9", x"03", x"03", x"ff", x"03", x"fd", x"fe",
    x"03", x"fd", x"fa", x"fc", x"fa", x"00", x"ff", x"01",
    x"ff", x"03", x"00", x"03", x"00", x"00", x"02", x"00",
    x"00", x"fb", x"fd", x"fb", x"fb", x"fe", x"02", x"ff",
    x"01", x"05", x"fe", x"fc", x"02", x"03", x"fa", x"01",
    x"fe", x"f7", x"f7", x"fc", x"fe", x"fd", x"fb", x"01",
    x"02", x"01", x"01", x"00", x"fc", x"fc", x"fb", x"00",
    x"fe", x"02", x"fc", x"02", x"fc", x"ff", x"fb", x"00",
    x"fe", x"05", x"02", x"fb", x"fc", x"00", x"fb", x"02",
    x"06", x"04", x"ff", x"fe", x"fe", x"03", x"ff", x"03",
    x"fc", x"f9", x"fe", x"fc", x"fb", x"03", x"fa", x"01",
    x"fc", x"fc", x"fc", x"03", x"04", x"fe", x"04", x"fd",
    x"fe", x"02", x"00", x"ff", x"fc", x"fc", x"fc", x"01",
    x"04", x"ff", x"f9", x"02", x"fe", x"f8", x"fe", x"fd",
    x"01", x"fe", x"04", x"ff", x"02", x"fd", x"fc", x"fd",
    x"fe", x"00", x"fd", x"01", x"fa", x"fc", x"fb", x"f9",
    x"fa", x"f5", x"ff", x"ff", x"fa", x"fa", x"fd", x"04",
    x"ff", x"f8", x"fd", x"fa", x"00", x"fd", x"03", x"02",
    x"01", x"fe", x"fc", x"00", x"fe", x"fb", x"fc", x"f9",
    x"00", x"fb", x"fe", x"fa", x"fc", x"00", x"fc", x"04",
    x"02", x"ff", x"f7", x"fd", x"fa", x"00", x"01", x"fe",
    x"fe", x"fa", x"00", x"00", x"fd", x"fc", x"01", x"fc",
    x"02", x"fb", x"fb", x"fb", x"01", x"f9", x"fa", x"fe",
    x"06", x"ff", x"fd", x"03", x"02", x"fc", x"04", x"00",
    x"ff", x"fe", x"fa", x"fa", x"ff", x"fb", x"03", x"ff",
    x"ff", x"f8", x"19", x"e9", x"e0", x"2a", x"bc", x"c0",
    x"05", x"d4", x"ea", x"fa", x"fa", x"c5", x"98", x"04",
    x"e8", x"f3", x"f5", x"e2", x"e8", x"d3", x"f2", x"fc",
    x"0e", x"25", x"31", x"bf", x"03", x"1f", x"21", x"10",
    x"df", x"18", x"0c", x"32", x"ff", x"1d", x"ff", x"ff",
    x"bb", x"c1", x"e2", x"ee", x"ce", x"fc", x"1e", x"27",
    x"34", x"0a", x"1e", x"ee", x"08", x"1d", x"27", x"fa",
    x"0a", x"3f", x"1d", x"28", x"54", x"57", x"1f", x"46",
    x"1d", x"d8", x"1b", x"0d", x"9a", x"d8", x"d2", x"e0",
    x"f3", x"e1", x"cc", x"e8", x"ca", x"67", x"8b", x"99",
    x"77", x"0a", x"f8", x"fc", x"c1", x"f4", x"0a", x"33",
    x"51", x"ea", x"c7", x"22", x"30", x"1d", x"27", x"2b",
    x"de", x"19", x"41", x"06", x"03", x"2d", x"25", x"4d",
    x"44", x"47", x"5f", x"21", x"11", x"db", x"db", x"3c",
    x"00", x"dd", x"fe", x"26", x"f7", x"e4", x"03", x"22",
    x"0a", x"12", x"3a", x"01", x"17", x"0e", x"09", x"f9",
    x"d6", x"2a", x"3f", x"1c", x"fa", x"0a", x"fe", x"f3",
    x"25", x"37", x"ea", x"0c", x"e8", x"e1", x"eb", x"df",
    x"3c", x"37", x"1e", x"fb", x"d2", x"cc", x"e1", x"e1",
    x"2a", x"05", x"01", x"fc", x"00", x"01", x"fd", x"fe",
    x"03", x"ff", x"d2", x"10", x"1b", x"f6", x"23", x"18",
    x"ee", x"f7", x"0d", x"ed", x"f2", x"f5", x"e5", x"be",
    x"ae", x"44", x"38", x"d0", x"e0", x"bf", x"1c", x"18",
    x"15", x"0b", x"0e", x"f5", x"05", x"02", x"25", x"06",
    x"01", x"d5", x"c6", x"12", x"7b", x"95", x"1e", x"27",
    x"15", x"3f", x"e6", x"e1", x"d4", x"d5", x"fa", x"fa",
    x"0f", x"ef", x"bd", x"c4", x"ed", x"e4", x"c5", x"a5",
    x"ec", x"eb", x"09", x"7f", x"fd", x"04", x"0a", x"d7",
    x"0a", x"db", x"c4", x"d7", x"b7", x"6c", x"d0", x"f8",
    x"d8", x"fa", x"22", x"f0", x"e6", x"a2", x"b1", x"ba",
    x"e5", x"ff", x"e7", x"f3", x"f5", x"f9", x"fa", x"f7",
    x"ff", x"fe", x"fb", x"01", x"20", x"16", x"2c", x"1c",
    x"39", x"46", x"e6", x"f5", x"c1", x"36", x"17", x"11",
    x"15", x"36", x"19", x"0f", x"ee", x"23", x"e5", x"f0",
    x"0f", x"2d", x"21", x"05", x"25", x"5b", x"24", x"1d",
    x"03", x"1b", x"0b", x"0e", x"ed", x"da", x"b3", x"74",
    x"d5", x"fb", x"2f", x"0b", x"10", x"38", x"39", x"41",
    x"52", x"dc", x"e4", x"ea", x"ea", x"0d", x"0b", x"0f",
    x"0b", x"10", x"d1", x"0a", x"14", x"26", x"1c", x"fc",
    x"1e", x"e4", x"e7", x"ed", x"ad", x"03", x"0a", x"d3",
    x"d2", x"ec", x"d9", x"b8", x"05", x"fd", x"f9", x"0c",
    x"00", x"06", x"f9", x"fb", x"fb", x"c4", x"15", x"30",
    x"10", x"f8", x"ec", x"0e", x"ef", x"f1", x"3d", x"21",
    x"1f", x"1d", x"29", x"06", x"1d", x"fc", x"ef", x"08",
    x"16", x"47", x"05", x"0a", x"1b", x"2d", x"1d", x"0f",
    x"fe", x"fb", x"fa", x"fd", x"fe", x"06", x"05", x"02",
    x"00", x"f9", x"f9", x"ee", x"c9", x"bf", x"e9", x"c2",
    x"87", x"a1", x"04", x"fe", x"02", x"eb", x"fe", x"e7",
    x"cd", x"ac", x"8f", x"09", x"0f", x"0c", x"c6", x"a3",
    x"92", x"e5", x"b7", x"b3", x"c2", x"08", x"1a", x"05",
    x"f6", x"f7", x"1f", x"0c", x"ff", x"fb", x"fd", x"c6",
    x"0d", x"f9", x"ec", x"96", x"a4", x"d5", x"d6", x"db",
    x"a4", x"c3", x"d7", x"f2", x"f0", x"08", x"0b", x"d2",
    x"d5", x"d3", x"f1", x"23", x"22", x"d7", x"1d", x"20",
    x"07", x"05", x"00", x"01", x"00", x"ff", x"ff", x"fb",
    x"04", x"00", x"03", x"03", x"02", x"fb", x"fc", x"01",
    x"ff", x"03", x"11", x"ea", x"f4", x"bd", x"c8", x"c1",
    x"92", x"c8", x"ef", x"37", x"1e", x"50", x"1b", x"21",
    x"2a", x"09", x"f7", x"e6", x"e1", x"fb", x"03", x"1f",
    x"30", x"2d", x"ca", x"00", x"33", x"2d", x"03", x"e7",
    x"0c", x"e4", x"df", x"e9", x"ed", x"df", x"3a", x"24",
    x"1f", x"b6", x"2a", x"2c", x"ec", x"01", x"18", x"17",
    x"af", x"c8", x"3d", x"2c", x"32", x"7b", x"3d", x"26",
    x"3f", x"30", x"40", x"05", x"1b", x"1e", x"01", x"2a",
    x"04", x"d4", x"fe", x"17", x"dd", x"cc", x"df", x"08",
    x"17", x"41", x"05", x"db", x"f3", x"11", x"27", x"1b",
    x"13", x"03", x"07", x"06", x"f9", x"f3", x"0f", x"08",
    x"1e", x"05", x"e5", x"06", x"e5", x"f4", x"e8", x"c6",
    x"df", x"23", x"0e", x"21", x"3a", x"1f", x"fd", x"fb",
    x"e3", x"e8", x"e4", x"20", x"e4", x"cc", x"0d", x"e3",
    x"da", x"24", x"cb", x"bc", x"f4", x"1e", x"fe", x"db",
    x"1e", x"2b", x"3b", x"26", x"0f", x"ee", x"cf", x"3a",
    x"00", x"0b", x"bb", x"e8", x"ef", x"c3", x"d6", x"f6",
    x"17", x"2e", x"f2", x"f4", x"16", x"ff", x"dd", x"33",
    x"f3", x"95", x"d9", x"0d", x"4a", x"c7", x"e5", x"fc",
    x"00", x"fa", x"fc", x"d3", x"f7", x"fc", x"e5", x"cb",
    x"e7", x"e6", x"e6", x"ec", x"0b", x"05", x"0d", x"e6",
    x"df", x"c8", x"aa", x"e8", x"d7", x"17", x"0b", x"ef",
    x"c9", x"fb", x"ba", x"0e", x"88", x"a9", x"04", x"c8",
    x"ad", x"28", x"1d", x"34", x"1f", x"4d", x"4b", x"f2",
    x"f4", x"33", x"0c", x"16", x"dc", x"e4", x"f4", x"d9",
    x"1c", x"35", x"26", x"18", x"0d", x"11", x"9a", x"d2",
    x"1e", x"ee", x"0a", x"17", x"1e", x"20", x"41", x"4f",
    x"4d", x"61", x"22", x"37", x"12", x"31", x"43", x"19",
    x"39", x"eb", x"1b", x"db", x"c8", x"d4", x"b6", x"cd",
    x"0c", x"fc", x"29", x"18", x"c6", x"c5", x"02", x"dc",
    x"c3", x"d7", x"ad", x"8d", x"c5", x"17", x"0c", x"9d",
    x"ee", x"0b", x"f7", x"f5", x"17", x"00", x"1d", x"0b",
    x"29", x"13", x"1b", x"fe", x"29", x"22", x"3b", x"a2",
    x"76", x"99", x"e9", x"0d", x"e6", x"2b", x"23", x"fb",
    x"c4", x"fd", x"06", x"de", x"1a", x"f5", x"0c", x"c2",
    x"22", x"00", x"03", x"00", x"ff", x"01", x"03", x"01",
    x"01", x"fb", x"23", x"55", x"32", x"1c", x"1d", x"f7",
    x"ed", x"f2", x"e6", x"11", x"36", x"e8", x"0f", x"24",
    x"ef", x"30", x"49", x"12", x"18", x"ff", x"f5", x"00",
    x"e4", x"b4", x"2b", x"30", x"e2", x"46", x"fb", x"01",
    x"1f", x"14", x"0c", x"b8", x"c5", x"05", x"21", x"0e",
    x"dc", x"11", x"f5", x"b8", x"08", x"ac", x"cb", x"ff",
    x"e5", x"f1", x"eb", x"eb", x"f1", x"cf", x"c5", x"cd",
    x"4b", x"09", x"14", x"37", x"f4", x"04", x"b4", x"f0",
    x"15", x"24", x"16", x"1d", x"0f", x"e9", x"f3", x"39",
    x"fe", x"bd", x"2b", x"32", x"2a", x"01", x"26", x"37",
    x"c5", x"be", x"b8", x"04", x"fe", x"02", x"00", x"fb",
    x"02", x"02", x"fe", x"fb", x"11", x"e7", x"ce", x"0d",
    x"d3", x"bc", x"e7", x"ed", x"c1", x"40", x"17", x"e1",
    x"2f", x"d2", x"be", x"74", x"3c", x"0c", x"23", x"f5",
    x"ed", x"27", x"45", x"3d", x"35", x"43", x"53", x"e8",
    x"f4", x"0f", x"0c", x"fb", x"e3", x"f7", x"e5", x"b7",
    x"f6", x"ea", x"fd", x"13", x"e4", x"e8", x"f5", x"cf",
    x"11", x"23", x"2f", x"17", x"19", x"03", x"4d", x"23",
    x"e2", x"b8", x"f8", x"c5", x"f9", x"b3", x"a0", x"cf",
    x"41", x"f1", x"c4", x"26", x"09", x"04", x"20", x"09",
    x"1a", x"ca", x"15", x"1f", x"fe", x"09", x"05", x"02",
    x"04", x"04", x"fc", x"fb", x"06", x"44", x"2e", x"2b",
    x"22", x"1e", x"18", x"17", x"18", x"f9", x"33", x"14",
    x"fe", x"fd", x"fb", x"f1", x"ef", x"0e", x"27", x"16",
    x"f1", x"1d", x"f1", x"fd", x"07", x"25", x"1c", x"35",
    x"09", x"ff", x"02", x"02", x"fd", x"04", x"03", x"fc",
    x"fd", x"1c", x"05", x"02", x"42", x"17", x"26", x"59",
    x"4a", x"28", x"25", x"1c", x"27", x"18", x"ff", x"03",
    x"19", x"fb", x"fb", x"0b", x"01", x"1a", x"15", x"1a",
    x"1f", x"3f", x"21", x"1f", x"eb", x"19", x"ba", x"14",
    x"f8", x"ef", x"ef", x"d5", x"d2", x"01", x"fc", x"0f",
    x"06", x"13", x"22", x"d1", x"d8", x"02", x"4f", x"23",
    x"d9", x"07", x"0b", x"d9", x"ec", x"f8", x"ce", x"4c",
    x"39", x"2a", x"09", x"18", x"e5", x"07", x"11", x"f4",
    x"09", x"02", x"03", x"05", x"01", x"05", x"03", x"06",
    x"06", x"05", x"02", x"f8", x"fe", x"01", x"04", x"fa",
    x"fc", x"ff", x"31", x"0a", x"2d", x"c0", x"f2", x"08",
    x"6d", x"b3", x"f4", x"08", x"32", x"18", x"23", x"18",
    x"2a", x"0e", x"0e", x"69", x"0b", x"38", x"17", x"ec",
    x"00", x"21", x"12", x"f3", x"f7", x"04", x"e6", x"f5",
    x"e8", x"c5", x"d2", x"d5", x"f9", x"f4", x"ee", x"e5",
    x"a9", x"f6", x"e8", x"f7", x"e4", x"dd", x"de", x"d3",
    x"0a", x"13", x"fb", x"fe", x"e0", x"48", x"34", x"28",
    x"07", x"e8", x"f0", x"d2", x"a8", x"f7", x"d0", x"fa",
    x"f6", x"22", x"16", x"e4", x"22", x"47", x"e8", x"02",
    x"34", x"d9", x"fd", x"f2", x"0a", x"06", x"df", x"d9",
    x"02", x"40", x"07", x"06", x"06", x"0b", x"d3", x"d1",
    x"e4", x"9f", x"42", x"4e", x"18", x"f8", x"21", x"13",
    x"e3", x"2b", x"d2", x"d4", x"ee", x"13", x"53", x"f2",
    x"e5", x"2d", x"ca", x"1b", x"22", x"f1", x"e4", x"13",
    x"31", x"f7", x"00", x"0e", x"dd", x"ab", x"ee", x"ae",
    x"e5", x"ec", x"03", x"bc", x"7d", x"fd", x"ad", x"a6",
    x"94", x"de", x"15", x"e6", x"f2", x"4c", x"fb", x"e0",
    x"0f", x"2c", x"08", x"f1", x"d5", x"d2", x"ea", x"84",
    x"31", x"00", x"e3", x"ef", x"d1", x"f1", x"40", x"4f",
    x"b9", x"b2", x"af", x"17", x"1c", x"f0", x"14", x"d1",
    x"ed", x"c2", x"27", x"20", x"40", x"0b", x"f4", x"15",
    x"27", x"fa", x"c3", x"d9", x"fb", x"1a", x"36", x"1e",
    x"e3", x"1e", x"38", x"e5", x"e2", x"b9", x"ea", x"d0",
    x"0b", x"23", x"0e", x"e0", x"69", x"e7", x"cc", x"f9",
    x"c0", x"da", x"65", x"af", x"41", x"11", x"03", x"32",
    x"0f", x"cb", x"e1", x"05", x"de", x"ee", x"01", x"0e",
    x"1c", x"fb", x"15", x"fa", x"97", x"ad", x"03", x"45",
    x"52", x"36", x"30", x"03", x"08", x"13", x"14", x"1a",
    x"39", x"ee", x"db", x"c8", x"e1", x"29", x"d8", x"bc",
    x"f2", x"7e", x"ea", x"cd", x"41", x"0f", x"d9", x"de",
    x"a6", x"c4", x"d7", x"ec", x"f6", x"9a", x"cf", x"c8",
    x"04", x"ff", x"0b", x"09", x"f8", x"3b", x"ff", x"16",
    x"26", x"d5", x"31", x"13", x"e4", x"d2", x"b1", x"1f",
    x"d8", x"f1", x"d6", x"b2", x"d6", x"19", x"3c", x"32",
    x"e2", x"d7", x"ae", x"01", x"0e", x"2f", x"18", x"30",
    x"2a", x"04", x"00", x"02", x"05", x"02", x"fe", x"04",
    x"05", x"ff", x"c9", x"db", x"a2", x"31", x"f0", x"20",
    x"cb", x"c9", x"b6", x"e8", x"08", x"1a", x"19", x"ed",
    x"10", x"ef", x"df", x"02", x"e7", x"e0", x"09", x"d6",
    x"be", x"f4", x"14", x"37", x"5c", x"f4", x"ff", x"d5",
    x"25", x"08", x"f4", x"da", x"d1", x"c8", x"01", x"cb",
    x"d9", x"07", x"03", x"20", x"d4", x"d6", x"c9", x"1e",
    x"fd", x"b8", x"e5", x"e0", x"e9", x"f0", x"ea", x"ef",
    x"02", x"64", x"c7", x"c3", x"25", x"1c", x"68", x"3d",
    x"10", x"de", x"13", x"38", x"0d", x"04", x"02", x"4c",
    x"3f", x"3d", x"f5", x"1c", x"0c", x"25", x"29", x"0f",
    x"f1", x"b0", x"c1", x"01", x"fa", x"fc", x"06", x"03",
    x"fe", x"fe", x"06", x"00", x"09", x"a2", x"a3", x"dd",
    x"e7", x"e3", x"f6", x"0c", x"f5", x"e6", x"d7", x"b6",
    x"00", x"d9", x"eb", x"ca", x"84", x"c2", x"d4", x"02",
    x"31", x"1a", x"00", x"26", x"29", x"42", x"33", x"20",
    x"a2", x"76", x"a9", x"82", x"bf", x"e3", x"00", x"05",
    x"dd", x"b1", x"bf", x"af", x"1d", x"0d", x"ed", x"f1",
    x"f9", x"1c", x"f8", x"1e", x"ae", x"db", x"df", x"59",
    x"39", x"15", x"52", x"f6", x"f2", x"ed", x"f4", x"f6",
    x"e6", x"06", x"18", x"d9", x"a1", x"9b", x"e3", x"dd",
    x"01", x"e1", x"15", x"05", x"f7", x"fc", x"fb", x"fc",
    x"fb", x"0a", x"f7", x"fd", x"00", x"f0", x"e5", x"d6",
    x"09", x"1b", x"01", x"04", x"01", x"0f", x"f2", x"1d",
    x"de", x"d9", x"d4", x"e9", x"1b", x"fd", x"0e", x"07",
    x"12", x"25", x"18", x"0a", x"f4", x"26", x"f8", x"eb",
    x"02", x"01", x"01", x"01", x"fb", x"03", x"03", x"fd",
    x"fb", x"f4", x"d1", x"c8", x"33", x"38", x"28", x"03",
    x"08", x"04", x"19", x"de", x"e5", x"fd", x"f5", x"0d",
    x"f4", x"ef", x"f8", x"e2", x"f1", x"09", x"0c", x"d6",
    x"da", x"34", x"42", x"3b", x"f4", x"1c", x"be", x"10",
    x"0e", x"15", x"e8", x"ea", x"ec", x"d0", x"d0", x"f7",
    x"fb", x"e8", x"fa", x"2b", x"10", x"0b", x"a1", x"ce",
    x"7f", x"14", x"13", x"23", x"1b", x"0a", x"b7", x"da",
    x"c8", x"b6", x"2f", x"20", x"18", x"f7", x"f2", x"ea",
    x"06", x"fe", x"02", x"02", x"fc", x"05", x"04", x"ff",
    x"fb", x"fc", x"02", x"04", x"fa", x"fb", x"fd", x"ff",
    x"fc", x"ff", x"2a", x"3a", x"b7", x"23", x"16", x"05",
    x"d4", x"d7", x"a8", x"1a", x"f5", x"3b", x"2c", x"07",
    x"f0", x"e5", x"d9", x"05", x"c1", x"0a", x"00", x"10",
    x"f4", x"08", x"c6", x"b7", x"d5", x"d1", x"e6", x"ed",
    x"1c", x"2c", x"25", x"16", x"e7", x"ec", x"e6", x"e6",
    x"04", x"f4", x"c7", x"c7", x"b9", x"b4", x"f7", x"1b",
    x"a3", x"7f", x"d0", x"00", x"08", x"fb", x"ba", x"eb",
    x"dd", x"01", x"06", x"ce", x"ca", x"d7", x"e7", x"fe",
    x"ed", x"02", x"f9", x"1d", x"4e", x"21", x"ce", x"46",
    x"27", x"2a", x"e5", x"0f", x"cc", x"02", x"16", x"39",
    x"17", x"0d", x"19", x"1c", x"00", x"f6", x"18", x"12",
    x"0c", x"07", x"c8", x"d4", x"df", x"e7", x"cb", x"21",
    x"17", x"19", x"38", x"46", x"1f", x"f8", x"cf", x"17",
    x"10", x"13", x"04", x"21", x"11", x"46", x"1c", x"9e",
    x"76", x"01", x"29", x"24", x"fd", x"0a", x"12", x"33",
    x"dc", x"14", x"a3", x"ad", x"c1", x"d9", x"c6", x"b2",
    x"4b", x"1c", x"0d", x"f8", x"1c", x"2f", x"d8", x"03",
    x"1f", x"25", x"0f", x"10", x"aa", x"f3", x"05", x"f4",
    x"f2", x"f0", x"2a", x"1c", x"20", x"13", x"08", x"fd",
    x"0c", x"09", x"f2", x"d0", x"cb", x"e5", x"03", x"2d",
    x"c4", x"fe", x"13", x"de", x"ec", x"cf", x"0e", x"ca",
    x"ea", x"0b", x"ed", x"ed", x"21", x"36", x"1e", x"0a",
    x"11", x"fd", x"1d", x"92", x"ef", x"de", x"10", x"31",
    x"cd", x"24", x"fc", x"fd", x"29", x"07", x"13", x"09",
    x"16", x"62", x"d1", x"dc", x"c3", x"a8", x"8b", x"92",
    x"1d", x"eb", x"ea", x"e2", x"f0", x"f9", x"d2", x"2d",
    x"2a", x"24", x"f8", x"0e", x"32", x"22", x"14", x"30",
    x"4c", x"1c", x"34", x"ec", x"e3", x"94", x"03", x"ff",
    x"3d", x"12", x"23", x"25", x"32", x"d8", x"5b", x"d4",
    x"c9", x"7d", x"d8", x"d3", x"cf", x"2a", x"1a", x"07",
    x"0a", x"ec", x"f3", x"d8", x"05", x"18", x"12", x"a5",
    x"15", x"00", x"06", x"0b", x"22", x"30", x"3a", x"32",
    x"1e", x"f8", x"18", x"23", x"0d", x"27", x"0d", x"0b",
    x"2d", x"04", x"2d", x"12", x"f3", x"32", x"1c", x"dd",
    x"92", x"c5", x"f7", x"8c", x"92", x"15", x"ca", x"d6",
    x"00", x"ff", x"ff", x"04", x"04", x"02", x"05", x"02",
    x"04", x"ff", x"00", x"21", x"45", x"e6", x"0b", x"f2",
    x"e6", x"c7", x"db", x"05", x"0a", x"eb", x"ee", x"00",
    x"32", x"3a", x"37", x"4c", x"5c", x"3b", x"ef", x"c6",
    x"06", x"40", x"b1", x"ca", x"e6", x"f6", x"e0", x"fb",
    x"e9", x"ee", x"10", x"f1", x"eb", x"24", x"d8", x"cf",
    x"cb", x"ca", x"f4", x"f6", x"cf", x"d4", x"f9", x"09",
    x"d7", x"b1", x"f4", x"97", x"a1", x"b0", x"d5", x"d4",
    x"ba", x"28", x"0f", x"fe", x"26", x"16", x"ea", x"20",
    x"31", x"27", x"2f", x"0c", x"ee", x"16", x"2f", x"4d",
    x"1f", x"4d", x"0b", x"fb", x"16", x"04", x"f3", x"08",
    x"ee", x"f1", x"1e", x"0f", x"01", x"0b", x"0b", x"0b",
    x"05", x"0d", x"05", x"07", x"c9", x"df", x"b6", x"c1",
    x"96", x"ba", x"de", x"ea", x"e4", x"13", x"d8", x"0f",
    x"30", x"1e", x"ff", x"49", x"19", x"f8", x"56", x"33",
    x"16", x"2f", x"44", x"25", x"55", x"49", x"50", x"ae",
    x"9e", x"bc", x"b9", x"95", x"98", x"af", x"91", x"98",
    x"0e", x"14", x"00", x"01", x"07", x"0f", x"de", x"ed",
    x"04", x"11", x"14", x"fa", x"0b", x"1a", x"17", x"fa",
    x"1f", x"30", x"17", x"47", x"33", x"71", x"3e", x"0b",
    x"eb", x"1d", x"09", x"46", x"48", x"2a", x"06", x"ff",
    x"05", x"a6", x"2a", x"fe", x"ff", x"03", x"08", x"fe",
    x"01", x"fe", x"fb", x"f9", x"fe", x"4b", x"f0", x"e4",
    x"04", x"f3", x"f8", x"e8", x"ec", x"f5", x"0d", x"e0",
    x"eb", x"33", x"e7", x"fa", x"27", x"2b", x"12", x"f0",
    x"f1", x"e3", x"f5", x"1b", x"27", x"dd", x"1c", x"31",
    x"fc", x"fc", x"05", x"00", x"02", x"00", x"fe", x"03",
    x"03", x"65", x"28", x"18", x"40", x"31", x"20", x"61",
    x"1c", x"35", x"cf", x"9f", x"9a", x"b0", x"9c", x"8c",
    x"c6", x"b4", x"e5", x"10", x"f9", x"fa", x"3d", x"14",
    x"10", x"4c", x"2e", x"27", x"e2", x"ea", x"e4", x"0b",
    x"11", x"38", x"fc", x"17", x"1d", x"fa", x"c8", x"cd",
    x"e9", x"02", x"30", x"e1", x"ed", x"1c", x"1f", x"d7",
    x"2a", x"0e", x"e6", x"db", x"1d", x"00", x"12", x"29",
    x"54", x"57", x"2d", x"20", x"36", x"01", x"14", x"2e",
    x"07", x"fc", x"fb", x"fa", x"02", x"f9", x"f9", x"fc",
    x"f9", x"03", x"07", x"09", x"03", x"07", x"06", x"03",
    x"00", x"08", x"f1", x"16", x"49", x"b8", x"fa", x"13",
    x"bd", x"e5", x"e1", x"ef", x"03", x"02", x"fd", x"2e",
    x"2f", x"e0", x"f2", x"37", x"39", x"36", x"45", x"1c",
    x"0e", x"20", x"b2", x"e7", x"20", x"dc", x"f3", x"e4",
    x"d5", x"f5", x"f6", x"e9", x"b8", x"bd", x"0c", x"1c",
    x"1e", x"03", x"ee", x"fb", x"11", x"ff", x"df", x"40",
    x"30", x"0f", x"32", x"07", x"0c", x"18", x"07", x"05",
    x"56", x"1a", x"c4", x"3b", x"fd", x"94", x"09", x"22",
    x"1c", x"c9", x"dd", x"06", x"52", x"04", x"20", x"53",
    x"36", x"2f", x"54", x"2d", x"36", x"05", x"fd", x"00",
    x"49", x"01", x"ed", x"59", x"25", x"2a", x"50", x"37",
    x"1f", x"eb", x"f1", x"ad", x"1d", x"28", x"2a", x"c7",
    x"f6", x"0b", x"21", x"03", x"f4", x"cf", x"c3", x"d1",
    x"82", x"13", x"0f", x"f8", x"fc", x"bc", x"39", x"42",
    x"5e", x"1f", x"2a", x"07", x"c4", x"f8", x"07", x"2d",
    x"33", x"46", x"c1", x"fc", x"16", x"98", x"f7", x"ea",
    x"49", x"c6", x"c3", x"57", x"15", x"f8", x"2e", x"46",
    x"e3", x"b7", x"19", x"02", x"04", x"28", x"10", x"03",
    x"23", x"0c", x"e3", x"89", x"84", x"de", x"cc", x"7a",
    x"11", x"f7", x"d1", x"d6", x"e1", x"dd", x"99", x"a5",
    x"ea", x"eb", x"b2", x"26", x"08", x"cd", x"04", x"0e",
    x"06", x"d6", x"29", x"35", x"a8", x"e2", x"1a", x"f8",
    x"df", x"c6", x"f5", x"d3", x"d3", x"f2", x"2c", x"00",
    x"21", x"16", x"eb", x"ff", x"b9", x"ce", x"c1", x"ed",
    x"24", x"6e", x"d3", x"f1", x"9b", x"f6", x"e9", x"db",
    x"f7", x"e7", x"eb", x"f6", x"f4", x"0e", x"09", x"f1",
    x"e5", x"e6", x"00", x"34", x"ca", x"f4", x"15", x"c2",
    x"ec", x"54", x"c5", x"bf", x"fe", x"09", x"e1", x"f5",
    x"45", x"27", x"06", x"4e", x"02", x"9f", x"3f", x"fb",
    x"de", x"17", x"ce", x"f9", x"37", x"25", x"2c", x"43",
    x"0e", x"15", x"4a", x"07", x"f8", x"b6", x"aa", x"a7",
    x"f3", x"b0", x"ab", x"3d", x"e8", x"0d", x"44", x"0f",
    x"08", x"0a", x"eb", x"eb", x"05", x"e1", x"e4", x"e0",
    x"ee", x"d4", x"04", x"1a", x"f8", x"f4", x"0b", x"10",
    x"31", x"14", x"76", x"12", x"f8", x"37", x"d5", x"fc",
    x"4e", x"ff", x"03", x"02", x"fe", x"03", x"05", x"ff",
    x"fd", x"ff", x"16", x"00", x"4c", x"d5", x"ea", x"e1",
    x"ff", x"ff", x"df", x"fa", x"cc", x"31", x"e7", x"10",
    x"2e", x"c2", x"0e", x"0f", x"f8", x"ce", x"25", x"f0",
    x"a1", x"cf", x"02", x"bf", x"d8", x"ea", x"28", x"03",
    x"f2", x"00", x"e5", x"de", x"e5", x"e0", x"0a", x"f3",
    x"47", x"e6", x"f9", x"58", x"e5", x"0e", x"23", x"f5",
    x"e4", x"f4", x"0e", x"f5", x"f8", x"2e", x"4d", x"e7",
    x"49", x"e0", x"d9", x"38", x"02", x"0a", x"df", x"e9",
    x"1f", x"05", x"d6", x"ec", x"41", x"03", x"19", x"23",
    x"07", x"ef", x"e6", x"f2", x"12", x"f8", x"05", x"00",
    x"e9", x"e7", x"ee", x"f6", x"f8", x"f4", x"fb", x"f6",
    x"fd", x"f5", x"f9", x"f6", x"f3", x"0d", x"15", x"eb",
    x"22", x"fe", x"07", x"18", x"15", x"10", x"39", x"65",
    x"02", x"33", x"72", x"f0", x"28", x"3f", x"9d", x"f6",
    x"d7", x"d7", x"fc", x"e6", x"ca", x"c5", x"ea", x"26",
    x"16", x"20", x"13", x"03", x"fc", x"0b", x"f7", x"fe",
    x"64", x"d7", x"06", x"36", x"05", x"18", x"0f", x"df",
    x"c6", x"17", x"fc", x"26", x"08", x"15", x"22", x"cb",
    x"04", x"1e", x"4d", x"37", x"e6", x"40", x"3c", x"dd",
    x"18", x"34", x"26", x"3a", x"f8", x"e5", x"1c", x"0c",
    x"0d", x"ce", x"1e", x"1a", x"f9", x"01", x"04", x"fa",
    x"fa", x"fa", x"fc", x"f1", x"ff", x"ee", x"f1", x"da",
    x"e9", x"d5", x"d7", x"01", x"ce", x"e9", x"2b", x"ff",
    x"19", x"75", x"1b", x"ea", x"51", x"f6", x"ee", x"55",
    x"ca", x"f8", x"2d", x"e8", x"ea", x"e7", x"b8", x"9c",
    x"02", x"00", x"fc", x"ff", x"06", x"fb", x"fb", x"05",
    x"ff", x"cc", x"e4", x"c2", x"c2", x"f8", x"16", x"f4",
    x"eb", x"26", x"22", x"e6", x"ee", x"e1", x"19", x"12",
    x"d2", x"ef", x"1d", x"c8", x"e4", x"e9", x"d9", x"0e",
    x"01", x"2d", x"2c", x"14", x"d5", x"bb", x"b4", x"b9",
    x"c7", x"ec", x"f8", x"e5", x"f5", x"0b", x"f6", x"f9",
    x"0d", x"0d", x"41", x"12", x"ff", x"2b", x"08", x"9b",
    x"78", x"c7", x"19", x"3b", x"ea", x"fe", x"ef", x"e6",
    x"20", x"ff", x"02", x"04", x"0e", x"0c", x"e7", x"ac",
    x"02", x"02", x"00", x"ff", x"fc", x"ff", x"03", x"fe",
    x"fe", x"fa", x"01", x"fc", x"07", x"fa", x"00", x"fc",
    x"fe", x"01", x"24", x"28", x"08", x"49", x"2b", x"ea",
    x"4b", x"4c", x"bf", x"1b", x"dd", x"1e", x"08", x"b2",
    x"f1", x"16", x"8a", x"b0", x"c5", x"ea", x"0d", x"e5",
    x"d6", x"0a", x"e3", x"f1", x"06", x"10", x"2c", x"14",
    x"06", x"1c", x"0c", x"e4", x"31", x"ff", x"3f", x"28",
    x"00", x"c9", x"e3", x"2b", x"d4", x"03", x"ef", x"44",
    x"12", x"f0", x"28", x"f9", x"1e", x"be", x"e7", x"c3",
    x"30", x"0b", x"f7", x"08", x"0b", x"de", x"56", x"f2",
    x"ef", x"1f", x"48", x"fe", x"e0", x"18", x"28", x"10",
    x"13", x"4f", x"f9", x"02", x"d4", x"0d", x"29", x"d4",
    x"48", x"28", x"d8", x"13", x"3a", x"29", x"e7", x"1b",
    x"0e", x"e8", x"e0", x"ef", x"17", x"3b", x"2c", x"11",
    x"26", x"31", x"1d", x"20", x"33", x"ca", x"20", x"3e",
    x"01", x"11", x"f4", x"ec", x"0f", x"19", x"33", x"3c",
    x"41", x"0f", x"02", x"26", x"41", x"0e", x"05", x"30",
    x"6a", x"55", x"00", x"5c", x"44", x"f5", x"3e", x"fc",
    x"ed", x"e2", x"15", x"0d", x"0d", x"16", x"2e", x"4e",
    x"59", x"2f", x"03", x"dd", x"1c", x"f4", x"05", x"ff",
    x"16", x"25", x"20", x"0d", x"f9", x"2d", x"27", x"05",
    x"e7", x"f7", x"ee", x"d8", x"09", x"05", x"af", x"e9",
    x"22", x"e2", x"8f", x"d5", x"da", x"ce", x"f8", x"22",
    x"27", x"e3", x"12", x"0e", x"05", x"0c", x"0b", x"18",
    x"37", x"34", x"67", x"28", x"34", x"40", x"21", x"04",
    x"c8", x"40", x"3f", x"2c", x"19", x"ff", x"20", x"ca",
    x"9d", x"d5", x"fa", x"f7", x"1e", x"16", x"22", x"06",
    x"e7", x"c8", x"65", x"fe", x"fa", x"b9", x"0a", x"13",
    x"f5", x"05", x"08", x"fe", x"d4", x"a5", x"d4", x"9d",
    x"a9", x"e5", x"65", x"4f", x"15", x"6d", x"35", x"fd",
    x"36", x"08", x"c5", x"c0", x"0a", x"2c", x"d7", x"30",
    x"36", x"d6", x"ef", x"0d", x"e9", x"f0", x"e0", x"18",
    x"26", x"39", x"f0", x"18", x"1c", x"02", x"19", x"37",
    x"fc", x"05", x"48", x"df", x"d5", x"42", x"fd", x"0c",
    x"34", x"c5", x"ca", x"e1", x"f9", x"b4", x"c3", x"1c",
    x"13", x"fc", x"d6", x"e6", x"08", x"b2", x"ea", x"27",
    x"df", x"fc", x"f1", x"0b", x"f8", x"14", x"f6", x"14",
    x"04", x"ff", x"01", x"fb", x"06", x"04", x"fb", x"02",
    x"fb", x"fb", x"16", x"0a", x"0f", x"fa", x"bc", x"f0",
    x"23", x"17", x"22", x"e5", x"10", x"34", x"fd", x"fb",
    x"0b", x"e4", x"d1", x"36", x"15", x"3d", x"4b", x"eb",
    x"fe", x"45", x"10", x"07", x"cf", x"fd", x"ff", x"2c",
    x"16", x"d9", x"f9", x"57", x"b6", x"96", x"10", x"13",
    x"19", x"fa", x"e9", x"f2", x"25", x"2f", x"12", x"fa",
    x"02", x"d5", x"1e", x"06", x"f0", x"e4", x"e3", x"e7",
    x"04", x"e9", x"0b", x"65", x"f6", x"e6", x"03", x"a6",
    x"bb", x"39", x"27", x"35", x"0a", x"0e", x"07", x"b5",
    x"cb", x"ab", x"26", x"fb", x"23", x"30", x"f6", x"f8",
    x"1e", x"17", x"1b", x"05", x"fe", x"05", x"f9", x"fe",
    x"fd", x"00", x"fb", x"09", x"f6", x"cf", x"b5", x"f0",
    x"d2", x"c4", x"f5", x"da", x"e9", x"1a", x"34", x"25",
    x"21", x"2a", x"1c", x"e2", x"d6", x"f7", x"16", x"ec",
    x"f1", x"df", x"cd", x"c0", x"7c", x"97", x"a9", x"ad",
    x"c6", x"c9", x"fd", x"ea", x"fe", x"1b", x"0a", x"16",
    x"df", x"d7", x"f8", x"02", x"fa", x"c8", x"02", x"10",
    x"55", x"07", x"f2", x"1a", x"12", x"e8", x"f8", x"05",
    x"02", x"28", x"d4", x"ee", x"0e", x"d0", x"de", x"19",
    x"bd", x"d8", x"ff", x"d1", x"fc", x"1e", x"35", x"16",
    x"0f", x"2d", x"dd", x"ca", x"03", x"02", x"fe", x"f9",
    x"fe", x"08", x"f4", x"09", x"f5", x"2c", x"6c", x"7a",
    x"34", x"4d", x"41", x"13", x"24", x"2b", x"68", x"36",
    x"17", x"05", x"07", x"08", x"14", x"f0", x"c7", x"1a",
    x"0f", x"2b", x"3c", x"2a", x"f1", x"05", x"ff", x"d8",
    x"ff", x"02", x"fd", x"fd", x"03", x"fc", x"fe", x"00",
    x"01", x"f9", x"06", x"ee", x"f8", x"36", x"46", x"df",
    x"dc", x"8d", x"fa", x"c6", x"ec", x"1c", x"d0", x"df",
    x"41", x"ee", x"a9", x"33", x"00", x"e5", x"1c", x"f0",
    x"dd", x"f9", x"5a", x"4f", x"06", x"3f", x"44", x"2d",
    x"21", x"3e", x"cf", x"f5", x"24", x"e8", x"03", x"0a",
    x"f2", x"e0", x"0e", x"f4", x"03", x"3a", x"30", x"c3",
    x"8b", x"05", x"0c", x"0e", x"00", x"13", x"28", x"1f",
    x"0c", x"22", x"27", x"12", x"2c", x"1c", x"33", x"22",
    x"fe", x"02", x"fa", x"08", x"02", x"04", x"fd", x"00",
    x"03", x"03", x"fe", x"fe", x"03", x"00", x"02", x"fe",
    x"08", x"03", x"01", x"07", x"12", x"f9", x"12", x"fc",
    x"c0", x"f2", x"06", x"f7", x"0e", x"3b", x"28", x"d3",
    x"b1", x"0c", x"d1", x"93", x"22", x"1c", x"21", x"40",
    x"43", x"56", x"1f", x"23", x"5c", x"ff", x"de", x"fb",
    x"23", x"f1", x"db", x"06", x"dd", x"00", x"1b", x"0f",
    x"fb", x"09", x"2e", x"25", x"28", x"fe", x"09", x"e0",
    x"af", x"eb", x"0e", x"10", x"f3", x"e5", x"14", x"2e",
    x"2e", x"25", x"1f", x"f3", x"01", x"fd", x"0e", x"0a",
    x"dc", x"f1", x"e6", x"b6", x"de", x"e9", x"c0", x"fc",
    x"cb", x"e7", x"2b", x"fc", x"f9", x"1a", x"31", x"40",
    x"00", x"4d", x"5a", x"da", x"d6", x"20", x"34", x"f8",
    x"fd", x"59", x"51", x"0c", x"04", x"eb", x"9b", x"18",
    x"fb", x"fd", x"d9", x"e2", x"f2", x"fa", x"cf", x"d5",
    x"ed", x"ed", x"f6", x"1a", x"fd", x"02", x"ff", x"b4",
    x"86", x"09", x"06", x"ed", x"25", x"30", x"14", x"e0",
    x"f0", x"01", x"12", x"f4", x"ef", x"ff", x"0b", x"11",
    x"da", x"cf", x"4d", x"f0", x"a1", x"27", x"0d", x"92",
    x"2d", x"03", x"0b", x"e3", x"41", x"fa", x"f1", x"16",
    x"01", x"f8", x"0a", x"15", x"26", x"d3", x"f7", x"fb",
    x"c4", x"05", x"08", x"fd", x"eb", x"fe", x"bc", x"f5",
    x"18", x"d5", x"e8", x"0f", x"f1", x"ed", x"04", x"e4",
    x"be", x"e0", x"ef", x"ad", x"e1", x"18", x"1a", x"11",
    x"0d", x"22", x"3b", x"02", x"11", x"41", x"e0", x"cb",
    x"f4", x"0c", x"13", x"21", x"11", x"5f", x"75", x"03",
    x"03", x"15", x"f8", x"16", x"dd", x"01", x"02", x"d7",
    x"d9", x"f1", x"d6", x"0b", x"de", x"bc", x"e9", x"af",
    x"cc", x"28", x"fd", x"1f", x"15", x"23", x"22", x"45",
    x"2f", x"34", x"59", x"13", x"30", x"52", x"fa", x"37",
    x"37", x"07", x"55", x"c5", x"fd", x"33", x"14", x"21",
    x"52", x"0e", x"2e", x"32", x"01", x"be", x"c9", x"0d",
    x"fa", x"f2", x"fd", x"c8", x"0a", x"25", x"40", x"87",
    x"00", x"35", x"74", x"11", x"f7", x"1e", x"e8", x"bf",
    x"e6", x"c3", x"f7", x"10", x"e9", x"25", x"f3", x"ab",
    x"ec", x"ee", x"a4", x"2e", x"07", x"eb", x"51", x"0c",
    x"20", x"0b", x"06", x"15", x"0e", x"01", x"15", x"f7",
    x"26", x"ff", x"05", x"fd", x"ff", x"00", x"03", x"02",
    x"00", x"00", x"2b", x"95", x"3f", x"42", x"35", x"3d",
    x"12", x"39", x"15", x"01", x"06", x"04", x"fb", x"0d",
    x"14", x"25", x"f6", x"14", x"cd", x"0f", x"59", x"d0",
    x"12", x"53", x"f4", x"13", x"33", x"11", x"27", x"fe",
    x"3c", x"1d", x"b8", x"5a", x"0e", x"d1", x"07", x"0c",
    x"35", x"0e", x"f0", x"c1", x"ec", x"d1", x"0f", x"e1",
    x"01", x"db", x"0a", x"01", x"aa", x"00", x"c9", x"99",
    x"f4", x"8d", x"05", x"4f", x"d4", x"e7", x"51", x"da",
    x"f5", x"0f", x"eb", x"25", x"1e", x"08", x"d7", x"f9",
    x"cf", x"db", x"0f", x"02", x"09", x"f8", x"e4", x"ca",
    x"3a", x"f6", x"f4", x"ff", x"01", x"06", x"05", x"ff",
    x"02", x"fb", x"02", x"06", x"1f", x"14", x"1b", x"df",
    x"fe", x"f9", x"ed", x"fd", x"f6", x"0d", x"08", x"12",
    x"1f", x"04", x"0d", x"13", x"f7", x"21", x"1f", x"34",
    x"25", x"d1", x"30", x"33", x"fc", x"4a", x"3c", x"e4",
    x"ea", x"e9", x"fd", x"18", x"f7", x"09", x"25", x"cd",
    x"db", x"eb", x"48", x"e9", x"00", x"09", x"f5", x"05",
    x"2c", x"02", x"16", x"fa", x"21", x"1d", x"31", x"1b",
    x"e3", x"19", x"cf", x"f3", x"07", x"e6", x"07", x"f7",
    x"fb", x"ea", x"45", x"09", x"f8", x"eb", x"4c", x"19",
    x"ee", x"41", x"19", x"f7", x"0a", x"12", x"13", x"12",
    x"0f", x"12", x"13", x"07", x"0d", x"3f", x"58", x"61",
    x"12", x"47", x"28", x"07", x"3b", x"29", x"49", x"03",
    x"fe", x"b3", x"0f", x"3d", x"ee", x"f2", x"0f", x"b9",
    x"02", x"24", x"98", x"e1", x"f8", x"96", x"08", x"4d",
    x"02", x"04", x"01", x"01", x"00", x"fc", x"fd", x"05",
    x"01", x"8f", x"0b", x"f8", x"35", x"ff", x"12", x"1f",
    x"05", x"0b", x"d5", x"fb", x"f1", x"3f", x"cc", x"e0",
    x"4e", x"d5", x"a4", x"29", x"f7", x"f8", x"5e", x"f8",
    x"01", x"08", x"fe", x"e4", x"40", x"15", x"49", x"ea",
    x"28", x"3a", x"49", x"19", x"15", x"0d", x"f1", x"db",
    x"01", x"ed", x"f3", x"01", x"de", x"28", x"5a", x"eb",
    x"8e", x"2e", x"ec", x"bb", x"1c", x"0a", x"fb", x"19",
    x"e9", x"e7", x"28", x"0b", x"2e", x"38", x"03", x"01",
    x"fd", x"05", x"05", x"04", x"06", x"03", x"06", x"03",
    x"00", x"01", x"fc", x"01", x"06", x"00", x"fa", x"02",
    x"f8", x"01", x"dc", x"fe", x"f3", x"be", x"cb", x"c1",
    x"98", x"8c", x"d9", x"d3", x"0f", x"94", x"fb", x"0b",
    x"58", x"0f", x"3b", x"56", x"00", x"1b", x"f1", x"06",
    x"17", x"0d", x"13", x"f6", x"dd", x"e7", x"05", x"fc",
    x"25", x"f5", x"ee", x"03", x"e2", x"ef", x"f1", x"fa",
    x"ec", x"2d", x"e0", x"1d", x"29", x"1d", x"0b", x"eb",
    x"93", x"c7", x"10", x"e5", x"f2", x"13", x"1c", x"10",
    x"01", x"e5", x"4d", x"ff", x"e1", x"20", x"d9", x"fa",
    x"2a", x"39", x"15", x"12", x"21", x"02", x"eb", x"08",
    x"fb", x"fa", x"fd", x"19", x"21", x"11", x"27", x"0c",
    x"24", x"13", x"14", x"3f", x"e2", x"f3", x"2d", x"2c",
    x"09", x"0d", x"40", x"1f", x"10", x"18", x"fb", x"38",
    x"e6", x"d7", x"26", x"f5", x"00", x"e0", x"0b", x"f3",
    x"2d", x"10", x"ce", x"25", x"eb", x"cf", x"08", x"df",
    x"00", x"ff", x"14", x"f2", x"16", x"09", x"05", x"e1",
    x"ed", x"e1", x"ed", x"0a", x"06", x"13", x"06", x"f4",
    x"26", x"1f", x"1e", x"1c", x"12", x"26", x"28", x"43",
    x"2b", x"0c", x"fa", x"00", x"0e", x"f2", x"ff", x"3e",
    x"e6", x"14", x"f9", x"d7", x"fa", x"ff", x"e7", x"0a",
    x"ce", x"ad", x"bf", x"d2", x"e2", x"1b", x"07", x"e3",
    x"32", x"21", x"04", x"21", x"f8", x"28", x"4a", x"01",
    x"2e", x"1d", x"36", x"fb", x"11", x"fb", x"16", x"07",
    x"0a", x"ea", x"86", x"ce", x"da", x"7d", x"da", x"e8",
    x"ec", x"1f", x"12", x"f2", x"ba", x"e9", x"f2", x"39",
    x"1e", x"ea", x"13", x"19", x"23", x"0a", x"0e", x"f6",
    x"0a", x"07", x"0b", x"e2", x"e8", x"fc", x"d8", x"06",
    x"ea", x"de", x"04", x"f1", x"be", x"03", x"16", x"f3",
    x"14", x"c9", x"40", x"51", x"47", x"fe", x"76", x"59",
    x"36", x"a9", x"ed", x"80", x"b7", x"eb", x"9d", x"1a",
    x"28", x"c2", x"1f", x"32", x"f0", x"f0", x"e6", x"55",
    x"2b", x"06", x"07", x"08", x"be", x"f7", x"c0", x"f2",
    x"c7", x"c0", x"d6", x"f4", x"db", x"d7", x"3d", x"11",
    x"e5", x"d6", x"f3", x"e5", x"e3", x"e9", x"e5", x"20",
    x"f5", x"ff", x"10", x"11", x"fb", x"b6", x"d8", x"22",
    x"1a", x"0a", x"e3", x"d5", x"d0", x"ae", x"ee", x"e3",
    x"fd", x"04", x"00", x"fc", x"fc", x"ff", x"fd", x"03",
    x"01", x"fe", x"3d", x"f3", x"f0", x"ca", x"f2", x"f2",
    x"e9", x"d2", x"f2", x"0e", x"0b", x"10", x"a1", x"91",
    x"af", x"0c", x"eb", x"e9", x"a5", x"f1", x"10", x"20",
    x"fd", x"da", x"04", x"fa", x"06", x"14", x"28", x"3b",
    x"ff", x"00", x"fa", x"9b", x"79", x"7b", x"1c", x"09",
    x"f7", x"2a", x"36", x"27", x"2b", x"16", x"e2", x"d4",
    x"4e", x"3d", x"fe", x"44", x"5c", x"26", x"09", x"30",
    x"bd", x"de", x"05", x"4a", x"19", x"14", x"08", x"ff",
    x"ed", x"ff", x"10", x"4e", x"e1", x"fe", x"05", x"cf",
    x"f6", x"dc", x"38", x"2a", x"3a", x"4a", x"a4", x"b2",
    x"99", x"56", x"6f", x"01", x"00", x"03", x"fd", x"f8",
    x"fe", x"f7", x"f6", x"01", x"14", x"04", x"1b", x"06",
    x"15", x"0e", x"26", x"30", x"07", x"3c", x"31", x"58",
    x"e2", x"4b", x"59", x"f4", x"f7", x"03", x"e0", x"bb",
    x"e1", x"d5", x"d6", x"ed", x"d7", x"f4", x"00", x"1c",
    x"0e", x"13", x"2b", x"0d", x"29", x"13", x"f8", x"0f",
    x"bc", x"f4", x"f2", x"0c", x"f5", x"13", x"15", x"01",
    x"0a", x"ca", x"f4", x"18", x"da", x"d8", x"27", x"ed",
    x"25", x"0e", x"a4", x"ab", x"df", x"f8", x"d3", x"c0",
    x"0d", x"ff", x"de", x"ff", x"f1", x"ed", x"17", x"07",
    x"01", x"f3", x"f1", x"e7", x"0b", x"02", x"f9", x"0a",
    x"fd", x"fc", x"fd", x"f8", x"ff", x"d8", x"f3", x"3b",
    x"fb", x"0b", x"12", x"ea", x"ca", x"0e", x"55", x"18",
    x"43", x"1f", x"2b", x"1b", x"4c", x"16", x"08", x"11",
    x"1e", x"13", x"3f", x"19", x"0c", x"0c", x"0c", x"27",
    x"fc", x"04", x"03", x"02", x"fd", x"04", x"02", x"fa",
    x"ff", x"e7", x"fe", x"0f", x"87", x"d8", x"e6", x"57",
    x"b6", x"9e", x"fc", x"1f", x"36", x"e3", x"28", x"26",
    x"22", x"10", x"f3", x"0c", x"08", x"22", x"ee", x"05",
    x"01", x"08", x"e8", x"11", x"2c", x"17", x"1d", x"de",
    x"f1", x"fa", x"e1", x"cd", x"d0", x"34", x"60", x"58",
    x"23", x"00", x"d3", x"0c", x"21", x"c8", x"e1", x"f9",
    x"b8", x"82", x"cb", x"0b", x"df", x"fd", x"f4", x"08",
    x"d7", x"e2", x"e2", x"e9", x"a7", x"dd", x"b6", x"c2",
    x"04", x"09", x"fd", x"07", x"02", x"09", x"08", x"09",
    x"04", x"fe", x"ff", x"f9", x"07", x"fe", x"00", x"fe",
    x"ff", x"f7", x"f3", x"01", x"ea", x"3d", x"22", x"15",
    x"1f", x"21", x"4c", x"20", x"2f", x"3f", x"11", x"0b",
    x"e7", x"12", x"07", x"dc", x"c4", x"eb", x"ff", x"08",
    x"1c", x"eb", x"ce", x"ff", x"05", x"1d", x"fb", x"e1",
    x"05", x"e0", x"e3", x"e0", x"bc", x"ed", x"c4", x"d9",
    x"d4", x"ab", x"d8", x"bc", x"dd", x"fd", x"13", x"f8",
    x"e9", x"d3", x"50", x"05", x"1f", x"16", x"e4", x"32",
    x"16", x"15", x"24", x"2f", x"34", x"34", x"fd", x"f6",
    x"01", x"41", x"41", x"fc", x"09", x"0c", x"e8", x"f8",
    x"01", x"f1", x"10", x"df", x"c2", x"37", x"40", x"38",
    x"e0", x"44", x"3f", x"e1", x"ec", x"d5", x"c4", x"95",
    x"7c", x"cb", x"a3", x"af", x"10", x"d4", x"e8", x"2f",
    x"22", x"0c", x"1f", x"02", x"09", x"2d", x"e8", x"d7",
    x"df", x"f0", x"0a", x"ea", x"2f", x"02", x"0c", x"d8",
    x"c0", x"36", x"09", x"08", x"03", x"f1", x"cf", x"ec",
    x"d8", x"a6", x"20", x"14", x"f3", x"0d", x"03", x"df",
    x"00", x"fb", x"fb", x"00", x"fd", x"00", x"02", x"fc",
    x"02", x"ff", x"fc", x"fe", x"ff", x"fb", x"fc", x"00",
    x"f9", x"fe", x"04", x"01", x"fa", x"fa", x"f9", x"fa",
    x"fa", x"02", x"00", x"fb", x"fa", x"fc", x"f8", x"fd",
    x"ff", x"ff", x"fa", x"fe", x"fd", x"02", x"f9", x"fb",
    x"fe", x"f8", x"fe", x"f9", x"01", x"00", x"02", x"fa",
    x"01", x"fd", x"fb", x"02", x"fd", x"01", x"fc", x"fe",
    x"03", x"fa", x"03", x"00", x"01", x"ff", x"fb", x"ff",
    x"fc", x"00", x"fb", x"fb", x"04", x"02", x"fb", x"01",
    x"01", x"00", x"04", x"ff", x"01", x"03", x"fb", x"fe",
    x"fb", x"05", x"ff", x"fd", x"02", x"fc", x"fb", x"01",
    x"01", x"fb", x"04", x"fc", x"fc", x"00", x"fa", x"fe",
    x"03", x"fc", x"ff", x"fd", x"fc", x"00", x"ff", x"03",
    x"fd", x"04", x"07", x"08", x"fc", x"fe", x"f9", x"fb",
    x"03", x"02", x"02", x"04", x"fa", x"fd", x"f9", x"fa",
    x"04", x"01", x"f9", x"fc", x"ff", x"fd", x"fc", x"fb",
    x"ff", x"fc", x"fb", x"01", x"fa", x"02", x"fa", x"03",
    x"fa", x"fc", x"ff", x"00", x"01", x"fe", x"fa", x"01",
    x"03", x"fa", x"01", x"03", x"03", x"05", x"fe", x"fc",
    x"fb", x"fc", x"ff", x"fb", x"04", x"00", x"00", x"03",
    x"fe", x"02", x"fa", x"fc", x"fe", x"01", x"01", x"ff",
    x"fd", x"01", x"fa", x"fa", x"02", x"fe", x"02", x"01",
    x"fe", x"01", x"00", x"fd", x"02", x"ff", x"fd", x"02",
    x"fe", x"fb", x"fe", x"fe", x"03", x"03", x"fd", x"02",
    x"fe", x"fc", x"fc", x"fa", x"02", x"ff", x"03", x"01",
    x"04", x"fb", x"01", x"02", x"ff", x"fd", x"fa", x"fe",
    x"fe", x"fc", x"02", x"03", x"02", x"fb", x"00", x"fd",
    x"02", x"fa", x"00", x"f9", x"00", x"fd", x"02", x"fd",
    x"fe", x"ff", x"03", x"fa", x"fc", x"03", x"fe", x"fd",
    x"fb", x"ff", x"01", x"f9", x"02", x"fd", x"ff", x"02",
    x"ff", x"fb", x"01", x"01", x"05", x"fb", x"03", x"05",
    x"fc", x"fc", x"fe", x"fc", x"02", x"fc", x"01", x"fc",
    x"ff", x"02", x"00", x"fe", x"01", x"00", x"f9", x"fe",
    x"fd", x"fd", x"ff", x"ff", x"fc", x"fd", x"fc", x"03",
    x"05", x"02", x"fb", x"01", x"02", x"ff", x"f9", x"fb",
    x"ff", x"f9", x"01", x"fa", x"03", x"fb", x"01", x"fe",
    x"fb", x"02", x"02", x"f9", x"fc", x"02", x"00", x"ff",
    x"01", x"00", x"f8", x"fd", x"fe", x"fc", x"fc", x"04",
    x"fd", x"fe", x"01", x"02", x"03", x"00", x"01", x"fc",
    x"04", x"ff", x"fb", x"02", x"f9", x"00", x"04", x"02",
    x"03", x"fa", x"01", x"01", x"fc", x"fb", x"04", x"fb",
    x"fd", x"03", x"fd", x"03", x"fc", x"04", x"ff", x"fc",
    x"00", x"ff", x"fd", x"fa", x"fd", x"01", x"f8", x"fb",
    x"00", x"fa", x"fa", x"01", x"05", x"fc", x"fc", x"02",
    x"02", x"01", x"02", x"04", x"00", x"fe", x"fe", x"00",
    x"fe", x"fe", x"ff", x"04", x"fe", x"fc", x"04", x"04",
    x"05", x"03", x"ff", x"03", x"fe", x"fc", x"fc", x"fe",
    x"fb", x"01", x"01", x"03", x"f9", x"fe", x"01", x"fd",
    x"fc", x"02", x"fe", x"fc", x"fd", x"fd", x"03", x"02",
    x"01", x"fd", x"fe", x"02", x"01", x"fc", x"fe", x"03",
    x"ff", x"02", x"fa", x"00", x"00", x"04", x"fa", x"05",
    x"02", x"01", x"02", x"fb", x"fd", x"fc", x"ff", x"fe",
    x"02", x"fd", x"fc", x"fc", x"fe", x"fd", x"fe", x"fa",
    x"03", x"fd", x"ff", x"fa", x"fb", x"f8", x"fd", x"01",
    x"00", x"02", x"03", x"fb", x"fd", x"fc", x"fd", x"05",
    x"04", x"04", x"04", x"fc", x"fe", x"01", x"fc", x"02",
    x"00", x"01", x"fc", x"02", x"fb", x"04", x"fe", x"05",
    x"fb", x"f9", x"02", x"03", x"fd", x"01", x"fb", x"fa",
    x"02", x"00", x"fc", x"fd", x"ff", x"fa", x"02", x"01",
    x"fe", x"f8", x"fc", x"fc", x"fd", x"04", x"fa", x"fb",
    x"01", x"01", x"fb", x"f9", x"f9", x"ff", x"01", x"00",
    x"00", x"fe", x"fa", x"fb", x"01", x"fd", x"01", x"02",
    x"fb", x"fa", x"ff", x"04", x"04", x"04", x"fc", x"ff",
    x"04", x"fa", x"00", x"01", x"01", x"06", x"01", x"05",
    x"02", x"ff", x"fd", x"02", x"fc", x"00", x"fb", x"f9",
    x"03", x"fa", x"03", x"fe", x"05", x"fc", x"fe", x"02",
    x"fa", x"f9", x"02", x"00", x"fa", x"fb", x"fc", x"04",
    x"fc", x"03", x"01", x"fc", x"00", x"fa", x"fe", x"fa",
    x"ff", x"fd", x"03", x"fd", x"02", x"00", x"f8", x"fc",
    x"fb", x"01", x"ff", x"02", x"01", x"fe", x"00", x"fc",
    x"f9", x"fc", x"fc", x"fa", x"03", x"02", x"fd", x"03",
    x"fe", x"fd", x"fe", x"fe", x"00", x"03", x"f8", x"01",
    x"fd", x"f7", x"fc", x"ff", x"fe", x"fe", x"ff", x"f6",
    x"fe", x"fb", x"ff", x"03", x"01", x"ff", x"fd", x"03",
    x"fd", x"01", x"fe", x"fb", x"fe", x"fc", x"ff", x"fc",
    x"01", x"ff", x"ff", x"fd", x"fe", x"fa", x"f7", x"f7",
    x"01", x"f9", x"f6", x"f9", x"fd", x"f9", x"fc", x"fb",
    x"03", x"02", x"00", x"fc", x"fa", x"02", x"fd", x"ff",
    x"03", x"f6", x"fc", x"02", x"fb", x"fe", x"04", x"ff",
    x"fc", x"fe", x"fc", x"fc", x"03", x"fe", x"00", x"00",
    x"02", x"fb", x"fd", x"fb", x"fd", x"02", x"fa", x"fe",
    x"fe", x"fc", x"03", x"01", x"fe", x"fd", x"04", x"00",
    x"ff", x"fa", x"fd", x"00", x"fc", x"fd", x"fc", x"03",
    x"fa", x"fe", x"00", x"fb", x"00", x"02", x"ff", x"03",
    x"01", x"02", x"fc", x"fb", x"fb", x"f5", x"fa", x"ff",
    x"fa", x"ff", x"fc", x"fb", x"fd", x"04", x"fe", x"00",
    x"fd", x"fe", x"01", x"fb", x"f9", x"04", x"00", x"05",
    x"fb", x"f9", x"01", x"02", x"f8", x"00", x"01", x"fc",
    x"04", x"fd", x"f9", x"fe", x"04", x"02", x"fe", x"01",
    x"00", x"fc", x"fd", x"03", x"04", x"fe", x"fc", x"fe",
    x"02", x"f9", x"fc", x"ff", x"fa", x"fd", x"fd", x"02",
    x"fc", x"01", x"ff", x"fc", x"04", x"03", x"05", x"02",
    x"04", x"04", x"00", x"03", x"04", x"04", x"fa", x"fa",
    x"fb", x"f7", x"f9", x"ff", x"02", x"fb", x"fb", x"02",
    x"fc", x"fc", x"fb", x"fc", x"fd", x"ff", x"ff", x"ff",
    x"00", x"fc", x"fa", x"fe", x"03", x"fd", x"f9", x"fa",
    x"fa", x"fc", x"00", x"01", x"fd", x"f9", x"03", x"fd",
    x"fb", x"f8", x"fe", x"03", x"04", x"04", x"fa", x"ff",
    x"fd", x"fd", x"fc", x"fa", x"01", x"01", x"fd", x"fe",
    x"ff", x"01", x"02", x"ff", x"ff", x"fd", x"01", x"01",
    x"fe", x"02", x"fe", x"ff", x"fe", x"fb", x"03", x"fc",
    x"00", x"fc", x"fe", x"01", x"f9", x"01", x"fc", x"02",
    x"fd", x"f8", x"fa", x"03", x"fc", x"fb", x"fe", x"fe",
    x"03", x"02", x"fc", x"fe", x"ff", x"fd", x"fa", x"04",
    x"f9", x"fd", x"ff", x"fd", x"fc", x"fc", x"00", x"fa",
    x"02", x"03", x"fd", x"04", x"fd", x"fe", x"fc", x"fa",
    x"fe", x"00", x"fc", x"f8", x"04", x"01", x"03", x"00",
    x"fa", x"fe", x"00", x"fc", x"00", x"fc", x"03", x"fb",
    x"fe", x"fb", x"01", x"ff", x"fd", x"fd", x"00", x"02",
    x"fe", x"ff", x"fa", x"fb", x"fa", x"fa", x"fc", x"fb",
    x"fd", x"fc", x"f9", x"f8", x"fd", x"fd", x"02", x"f7",
    x"fa", x"fd", x"ff", x"fd", x"fe", x"fc", x"fe", x"fe",
    x"fc", x"fb", x"fc", x"01", x"ff", x"02", x"00", x"01",
    x"04", x"01", x"01", x"fa", x"02", x"03", x"f7", x"ff",
    x"fc", x"ff", x"ff", x"fc", x"02", x"01", x"f9", x"fc",
    x"fc", x"ff", x"fa", x"fa", x"fe", x"02", x"01", x"fc",
    x"01", x"fc", x"01", x"fc", x"f5", x"fb", x"fc", x"fb",
    x"04", x"02", x"02", x"03", x"fd", x"fc", x"02", x"00",
    x"00", x"03", x"ff", x"fe", x"03", x"ff", x"fb", x"02",
    x"04", x"fc", x"ff", x"02", x"02", x"fe", x"ff", x"fe",
    x"fc", x"01", x"f8", x"01", x"02", x"00", x"00", x"fd",
    x"fc", x"fe", x"fe", x"fc", x"fd", x"f9", x"00", x"ff",
    x"fb", x"f8", x"fc", x"f7", x"ff", x"fd", x"fc", x"01",
    x"fe", x"fd", x"01", x"04", x"00", x"fc", x"fa", x"05",
    x"03", x"00", x"fd", x"fb", x"04", x"00", x"f9", x"00",
    x"00", x"ff", x"fd", x"00", x"ff", x"03", x"ff", x"fc",
    x"05", x"05", x"fe", x"03", x"05", x"ff", x"ff", x"05",
    x"03", x"05", x"00", x"00", x"01", x"01", x"02", x"04",
    x"01", x"fe", x"fe", x"fd", x"f8", x"fd", x"fe", x"01",
    x"ff", x"04", x"ff", x"ff", x"fa", x"fa", x"02", x"04",
    x"ff", x"fb", x"fe", x"fb", x"02", x"fc", x"fc", x"ff",
    x"fc", x"ff", x"ff", x"04", x"01", x"fb", x"fb", x"fc",
    x"fd", x"fd", x"01", x"00", x"ff", x"01", x"00", x"fd",
    x"ff", x"fb", x"01", x"01", x"fc", x"fa", x"fa", x"fb",
    x"fc", x"fd", x"fa", x"fa", x"00", x"fa", x"03", x"fd",
    x"fe", x"f9", x"f9", x"f9", x"fc", x"fc", x"fc", x"00",
    x"fc", x"02", x"ff", x"fa", x"fa", x"fb", x"fd", x"fd",
    x"fd", x"fd", x"00", x"ff", x"fd", x"00", x"03", x"f9",
    x"fd", x"fa", x"f8", x"fb", x"ff", x"fe", x"00", x"01",
    x"ff", x"fd", x"01", x"00", x"fb", x"02", x"00", x"fb",
    x"fd", x"ff", x"00", x"01", x"fa", x"ff", x"00", x"fb",
    x"fa", x"03", x"fa", x"01", x"fd", x"fc", x"fb", x"ff",
    x"01", x"02", x"fc", x"fc", x"ff", x"fe", x"01", x"fb",
    x"fe", x"fc", x"ff", x"04", x"02", x"01", x"03", x"03",
    x"db", x"c8", x"12", x"d9", x"b5", x"2b", x"03", x"df",
    x"12", x"18", x"18", x"f4", x"12", x"d9", x"0d", x"fb",
    x"2a", x"53", x"28", x"1a", x"28", x"11", x"14", x"25",
    x"0a", x"15", x"0a", x"c5", x"05", x"f8", x"cf", x"fa",
    x"fb", x"00", x"db", x"b2", x"1d", x"24", x"21", x"34",
    x"36", x"3c", x"0d", x"38", x"3f", x"ec", x"a8", x"bf",
    x"1c", x"db", x"65", x"28", x"00", x"9c", x"ff", x"c0",
    x"ca", x"a6", x"bb", x"ef", x"f6", x"fe", x"0e", x"08",
    x"0a", x"0b", x"1f", x"20", x"05", x"30", x"25", x"17",
    x"0a", x"02", x"0c", x"1c", x"f6", x"e6", x"24", x"ff",
    x"f3", x"eb", x"e2", x"f7", x"ed", x"19", x"36", x"13",
    x"fb", x"21", x"e2", x"16", x"32", x"d2", x"30", x"37",
    x"57", x"23", x"eb", x"7b", x"d4", x"eb", x"be", x"da",
    x"0d", x"3a", x"19", x"3b", x"00", x"f2", x"fb", x"fa",
    x"f3", x"19", x"3e", x"24", x"33", x"1a", x"08", x"3c",
    x"0e", x"f9", x"1a", x"00", x"07", x"5b", x"0c", x"28",
    x"29", x"19", x"18", x"29", x"24", x"19", x"1d", x"f0",
    x"de", x"d9", x"fe", x"a2", x"be", x"06", x"c7", x"e3",
    x"f0", x"8f", x"73", x"de", x"a8", x"81", x"f9", x"10",
    x"06", x"fc", x"ff", x"fc", x"fe", x"fd", x"01", x"ff",
    x"00", x"03", x"2a", x"33", x"2c", x"09", x"e7", x"f0",
    x"f4", x"f4", x"f6", x"f0", x"0d", x"18", x"fe", x"e0",
    x"19", x"13", x"a2", x"b3", x"f0", x"e0", x"22", x"18",
    x"08", x"e6", x"45", x"3d", x"5d", x"04", x"10", x"f6",
    x"fb", x"ea", x"eb", x"e2", x"e1", x"e7", x"cf", x"83",
    x"a9", x"e5", x"90", x"9a", x"24", x"d9", x"e4", x"23",
    x"16", x"cf", x"2d", x"1b", x"f4", x"01", x"07", x"31",
    x"13", x"fe", x"0a", x"de", x"ef", x"fb", x"28", x"32",
    x"16", x"d7", x"04", x"12", x"e7", x"d2", x"d6", x"0b",
    x"ca", x"de", x"04", x"06", x"08", x"13", x"14", x"07",
    x"ea", x"0f", x"65", x"08", x"05", x"01", x"fe", x"01",
    x"00", x"05", x"ff", x"fa", x"37", x"5b", x"5c", x"4c",
    x"34", x"18", x"33", x"16", x"15", x"25", x"0a", x"19",
    x"f5", x"02", x"f3", x"d4", x"e0", x"c8", x"27", x"0a",
    x"24", x"1b", x"14", x"20", x"2a", x"19", x"26", x"4a",
    x"3a", x"26", x"28", x"27", x"23", x"1a", x"fc", x"18",
    x"ac", x"e2", x"10", x"c1", x"c2", x"f7", x"ea", x"e1",
    x"f9", x"dd", x"fb", x"f1", x"fb", x"db", x"aa", x"ff",
    x"09", x"33", x"d4", x"15", x"ff", x"d4", x"f3", x"f8",
    x"ec", x"e6", x"19", x"d1", x"21", x"36", x"15", x"0e",
    x"17", x"32", x"3d", x"0f", x"04", x"ff", x"fd", x"fb",
    x"f9", x"02", x"f7", x"fa", x"08", x"12", x"26", x"2e",
    x"09", x"03", x"14", x"15", x"25", x"26", x"f0", x"75",
    x"3f", x"15", x"13", x"11", x"25", x"ea", x"e0", x"16",
    x"05", x"5f", x"f2", x"ec", x"e0", x"bf", x"d3", x"f1",
    x"f8", x"01", x"05", x"ff", x"fb", x"fd", x"01", x"02",
    x"ff", x"de", x"31", x"23", x"f1", x"16", x"25", x"2b",
    x"d0", x"d2", x"de", x"f2", x"1e", x"dd", x"fc", x"0d",
    x"2f", x"10", x"ec", x"2e", x"4b", x"58", x"40", x"32",
    x"41", x"00", x"36", x"4c", x"26", x"e2", x"1e", x"0b",
    x"fd", x"0d", x"13", x"ea", x"f8", x"04", x"08", x"e5",
    x"1a", x"0e", x"22", x"1f", x"2b", x"4b", x"5e", x"f2",
    x"eb", x"2a", x"e1", x"83", x"f3", x"d2", x"aa", x"f5",
    x"f3", x"0d", x"e1", x"f7", x"0f", x"e2", x"f9", x"da",
    x"08", x"06", x"00", x"06", x"ff", x"fc", x"fd", x"08",
    x"fe", x"f7", x"f9", x"ff", x"02", x"fe", x"fd", x"ff",
    x"fd", x"fe", x"e6", x"d5", x"e0", x"02", x"fd", x"03",
    x"1e", x"f3", x"16", x"e3", x"f6", x"36", x"eb", x"0d",
    x"19", x"fa", x"1b", x"17", x"fb", x"f8", x"20", x"00",
    x"ec", x"ef", x"26", x"08", x"e9", x"10", x"17", x"13",
    x"0c", x"dd", x"1c", x"32", x"dd", x"0f", x"a8", x"78",
    x"8f", x"c6", x"bd", x"c4", x"f7", x"0d", x"f9", x"b7",
    x"cf", x"e8", x"e0", x"bc", x"e2", x"f7", x"1a", x"30",
    x"c3", x"b2", x"f4", x"f6", x"bd", x"ed", x"18", x"f2",
    x"09", x"30", x"1b", x"19", x"0c", x"34", x"2f", x"01",
    x"41", x"4f", x"b4", x"84", x"a8", x"e6", x"b0", x"de",
    x"0d", x"bd", x"ca", x"d9", x"d9", x"05", x"f9", x"15",
    x"02", x"22", x"10", x"06", x"c6", x"1c", x"d6", x"d9",
    x"22", x"09", x"11", x"08", x"05", x"66", x"30", x"13",
    x"08", x"20", x"27", x"94", x"48", x"35", x"f1", x"cb",
    x"f3", x"df", x"d1", x"e9", x"14", x"1b", x"29", x"ee",
    x"cb", x"de", x"07", x"c2", x"cf", x"2f", x"0a", x"17",
    x"40", x"08", x"a4", x"2d", x"38", x"f2", x"22", x"19",
    x"c7", x"ff", x"1b", x"26", x"ec", x"24", x"1b", x"db",
    x"08", x"0e", x"06", x"ce", x"b3", x"fc", x"01", x"e0",
    x"1c", x"ec", x"bf", x"fe", x"0b", x"e8", x"0d", x"d8",
    x"c9", x"17", x"30", x"17", x"0f", x"f9", x"04", x"00",
    x"ab", x"17", x"2d", x"15", x"2b", x"24", x"18", x"17",
    x"d2", x"da", x"0b", x"c8", x"cc", x"d5", x"f3", x"10",
    x"e9", x"eb", x"ed", x"e1", x"da", x"98", x"3a", x"2c",
    x"01", x"36", x"f9", x"f5", x"08", x"ee", x"e6", x"f0",
    x"f9", x"f8", x"25", x"03", x"2b", x"3c", x"06", x"32",
    x"09", x"e9", x"ee", x"0e", x"05", x"fd", x"02", x"ef",
    x"d5", x"85", x"0c", x"c9", x"c9", x"31", x"ea", x"a5",
    x"3f", x"12", x"cc", x"1c", x"14", x"fc", x"3a", x"14",
    x"d8", x"05", x"ef", x"be", x"3f", x"31", x"e5", x"e7",
    x"f4", x"ff", x"e8", x"01", x"04", x"ef", x"de", x"a8",
    x"f0", x"da", x"4d", x"2b", x"ef", x"3b", x"1c", x"d3",
    x"26", x"bf", x"b1", x"01", x"b9", x"cb", x"ac", x"1f",
    x"0e", x"03", x"1a", x"fc", x"ce", x"27", x"cd", x"8f",
    x"2e", x"11", x"2c", x"17", x"2b", x"42", x"1a", x"57",
    x"5e", x"fc", x"04", x"00", x"fa", x"04", x"04", x"04",
    x"04", x"00", x"26", x"89", x"d1", x"84", x"a7", x"d2",
    x"fb", x"e0", x"d5", x"f3", x"00", x"36", x"29", x"37",
    x"34", x"23", x"29", x"f2", x"05", x"01", x"d1", x"27",
    x"f1", x"d6", x"0f", x"ec", x"f7", x"bd", x"e8", x"17",
    x"d9", x"32", x"38", x"d4", x"15", x"1d", x"ec", x"13",
    x"0e", x"fb", x"fd", x"35", x"e4", x"45", x"3e", x"47",
    x"fb", x"f6", x"38", x"0b", x"29", x"5a", x"40", x"4f",
    x"46", x"12", x"f5", x"ec", x"0a", x"ce", x"be", x"1f",
    x"0f", x"b7", x"f5", x"c8", x"06", x"09", x"e4", x"20",
    x"28", x"5a", x"c4", x"ff", x"08", x"ed", x"30", x"05",
    x"e8", x"4c", x"28", x"01", x"01", x"fe", x"fc", x"fa",
    x"ff", x"fb", x"fc", x"fb", x"a9", x"c7", x"03", x"e7",
    x"d9", x"0c", x"0e", x"02", x"f4", x"31", x"1c", x"e5",
    x"0a", x"e5", x"0d", x"19", x"00", x"f4", x"b5", x"df",
    x"db", x"b2", x"e2", x"9a", x"bb", x"c6", x"df", x"00",
    x"04", x"2a", x"ff", x"ff", x"15", x"f5", x"de", x"ea",
    x"44", x"e8", x"9a", x"19", x"12", x"aa", x"fd", x"d2",
    x"c3", x"11", x"f4", x"0b", x"01", x"f5", x"18", x"0e",
    x"3a", x"ef", x"09", x"0c", x"e2", x"29", x"1a", x"d5",
    x"12", x"12", x"02", x"23", x"20", x"ee", x"07", x"0b",
    x"34", x"01", x"e6", x"23", x"06", x"fc", x"05", x"02",
    x"f9", x"fa", x"02", x"fc", x"06", x"03", x"a6", x"85",
    x"dd", x"f5", x"e8", x"ff", x"bf", x"d1", x"e6", x"f2",
    x"e0", x"0c", x"12", x"ff", x"d8", x"15", x"0e", x"cc",
    x"fc", x"0d", x"b7", x"0c", x"db", x"e2", x"8a", x"7e",
    x"05", x"ff", x"05", x"04", x"fb", x"01", x"fb", x"01",
    x"01", x"cf", x"d9", x"f9", x"e4", x"13", x"fe", x"0d",
    x"da", x"cc", x"3f", x"03", x"f8", x"f2", x"0d", x"16",
    x"e6", x"19", x"e5", x"1e", x"09", x"07", x"3b", x"0f",
    x"1b", x"3c", x"2d", x"14", x"fa", x"06", x"f3", x"02",
    x"05", x"e3", x"fa", x"e1", x"b7", x"06", x"31", x"2b",
    x"17", x"f4", x"24", x"fc", x"eb", x"3b", x"0f", x"df",
    x"1f", x"f3", x"fb", x"2b", x"0d", x"09", x"04", x"15",
    x"ec", x"1d", x"13", x"e0", x"16", x"0c", x"e4", x"ea",
    x"03", x"02", x"06", x"fb", x"07", x"03", x"00", x"ff",
    x"00", x"fb", x"05", x"00", x"03", x"01", x"02", x"fb",
    x"00", x"fd", x"00", x"fe", x"1b", x"2e", x"08", x"05",
    x"19", x"4d", x"66", x"ef", x"bf", x"eb", x"fb", x"d7",
    x"5b", x"e3", x"b6", x"5d", x"cb", x"f0", x"2a", x"e4",
    x"cb", x"ff", x"de", x"c1", x"c5", x"08", x"22", x"34",
    x"d3", x"0d", x"23", x"f2", x"15", x"18", x"26", x"1f",
    x"f1", x"d6", x"1c", x"e6", x"e5", x"ee", x"e1", x"69",
    x"40", x"01", x"1d", x"29", x"a6", x"cb", x"a3", x"9c",
    x"2c", x"0b", x"9a", x"fb", x"c9", x"da", x"05", x"f0",
    x"ec", x"fa", x"2a", x"4b", x"f6", x"33", x"3b", x"d7",
    x"47", x"5c", x"df", x"09", x"cf", x"1f", x"cb", x"ca",
    x"1c", x"c1", x"9c", x"2d", x"f8", x"d1", x"ea", x"ef",
    x"cd", x"d6", x"d2", x"c5", x"1b", x"20", x"1d", x"4b",
    x"2e", x"0e", x"0d", x"4b", x"fe", x"f5", x"19", x"16",
    x"14", x"00", x"03", x"f2", x"ff", x"c2", x"3b", x"f1",
    x"ce", x"f2", x"d1", x"cc", x"e8", x"0d", x"0c", x"f3",
    x"21", x"df", x"e8", x"e5", x"db", x"fd", x"0f", x"15",
    x"fd", x"f9", x"f9", x"fa", x"ff", x"f8", x"f9", x"fd",
    x"fa", x"fc", x"02", x"f9", x"fb", x"fd", x"fe", x"fa",
    x"ff", x"fc", x"fe", x"03", x"fb", x"fb", x"fc", x"fa",
    x"04", x"fc", x"fc", x"f6", x"fa", x"f9", x"fb", x"f4",
    x"ff", x"fc", x"f9", x"ff", x"03", x"01", x"fa", x"ff",
    x"fe", x"01", x"f9", x"fe", x"fd", x"fe", x"01", x"fa",
    x"fa", x"fc", x"fe", x"fc", x"03", x"fa", x"fd", x"f9",
    x"00", x"fb", x"02", x"fc", x"f8", x"fc", x"fb", x"01",
    x"fe", x"03", x"fb", x"02", x"fb", x"04", x"00", x"04",
    x"01", x"02", x"fe", x"fc", x"02", x"fc", x"03", x"fd",
    x"fd", x"ff", x"fc", x"fa", x"00", x"ff", x"fb", x"fe",
    x"fb", x"fe", x"fd", x"03", x"fd", x"ff", x"ff", x"fb",
    x"fa", x"02", x"fa", x"fa", x"fe", x"fa", x"00", x"01",
    x"fe", x"fb", x"fa", x"fe", x"fb", x"ff", x"fb", x"02",
    x"fc", x"fc", x"04", x"fc", x"f7", x"fe", x"fe", x"02",
    x"fc", x"fd", x"f8", x"ff", x"f9", x"02", x"fb", x"ff",
    x"f8", x"05", x"01", x"fb", x"fb", x"fb", x"00", x"fa",
    x"fc", x"fc", x"ff", x"ff", x"fd", x"fd", x"fb", x"01",
    x"01", x"fb", x"fa", x"ff", x"01", x"ff", x"fc", x"fe",
    x"ff", x"fb", x"01", x"ff", x"fc", x"04", x"05", x"00",
    x"ff", x"05", x"fc", x"ff", x"ff", x"fb", x"fe", x"04",
    x"fa", x"02", x"fe", x"fe", x"02", x"f8", x"02", x"01",
    x"ff", x"fd", x"f6", x"ff", x"fc", x"00", x"ff", x"ff",
    x"fd", x"fe", x"03", x"fb", x"fd", x"fe", x"00", x"01",
    x"03", x"00", x"fd", x"fc", x"fc", x"fd", x"fa", x"fc",
    x"fd", x"00", x"fd", x"ff", x"fd", x"ff", x"ff", x"fb",
    x"fb", x"fe", x"fe", x"fa", x"fd", x"fc", x"fd", x"fa",
    x"fe", x"fb", x"f9", x"fe", x"fa", x"fb", x"ff", x"fe",
    x"f9", x"f7", x"02", x"fc", x"01", x"fe", x"00", x"fd",
    x"fd", x"00", x"fe", x"00", x"f7", x"ff", x"f9", x"fb",
    x"ff", x"fa", x"00", x"05", x"01", x"03", x"fe", x"fc",
    x"fe", x"05", x"05", x"00", x"03", x"fd", x"fd", x"00",
    x"04", x"fe", x"04", x"fe", x"fc", x"ff", x"ff", x"fa",
    x"00", x"00", x"fb", x"fe", x"f7", x"f6", x"ff", x"05",
    x"f9", x"fb", x"fc", x"f9", x"04", x"fb", x"02", x"fd",
    x"00", x"03", x"fc", x"03", x"fb", x"fc", x"04", x"fa",
    x"fb", x"00", x"fa", x"ff", x"03", x"01", x"ff", x"00",
    x"ff", x"ff", x"fa", x"f4", x"02", x"fc", x"01", x"02",
    x"fe", x"fd", x"fc", x"fc", x"fa", x"f9", x"01", x"f9",
    x"fd", x"ff", x"fa", x"ff", x"fc", x"ff", x"ff", x"f7",
    x"01", x"02", x"01", x"fd", x"04", x"ff", x"03", x"fe",
    x"04", x"02", x"00", x"05", x"ff", x"03", x"fd", x"02",
    x"04", x"02", x"f8", x"fd", x"02", x"f7", x"fa", x"02",
    x"fd", x"fa", x"fd", x"fe", x"fe", x"fa", x"fc", x"fb",
    x"fd", x"fd", x"f6", x"01", x"f9", x"f6", x"03", x"fa",
    x"01", x"fe", x"01", x"00", x"01", x"04", x"02", x"fd",
    x"fe", x"fc", x"ff", x"fd", x"00", x"fe", x"fe", x"fc",
    x"fa", x"fa", x"fe", x"fc", x"f9", x"03", x"ff", x"00",
    x"fc", x"02", x"f9", x"02", x"fe", x"f9", x"04", x"fd",
    x"ff", x"01", x"fc", x"fb", x"01", x"fe", x"fb", x"fe",
    x"fb", x"03", x"fb", x"fc", x"fd", x"01", x"00", x"fe",
    x"03", x"ff", x"fd", x"fd", x"fe", x"00", x"fa", x"fe",
    x"fa", x"00", x"fc", x"ff", x"fe", x"fb", x"fb", x"ff",
    x"fe", x"01", x"02", x"fd", x"00", x"fa", x"fc", x"03",
    x"fc", x"00", x"03", x"fc", x"03", x"04", x"fc", x"fd",
    x"fe", x"03", x"fb", x"01", x"fc", x"01", x"00", x"fd",
    x"03", x"02", x"fe", x"fc", x"04", x"02", x"ff", x"f7",
    x"fe", x"05", x"01", x"01", x"fb", x"01", x"03", x"ff",
    x"fc", x"fb", x"fe", x"fc", x"fb", x"f6", x"fe", x"04",
    x"fb", x"ff", x"02", x"fb", x"fd", x"ff", x"f8", x"f9",
    x"fe", x"fc", x"00", x"f8", x"ff", x"ff", x"f9", x"fd",
    x"fc", x"00", x"ff", x"fe", x"ff", x"fc", x"f8", x"00",
    x"01", x"fe", x"fd", x"01", x"04", x"05", x"04", x"ff",
    x"fc", x"fe", x"fe", x"fc", x"f6", x"fd", x"fb", x"fd",
    x"00", x"fc", x"fc", x"f7", x"fc", x"00", x"01", x"fb",
    x"fb", x"fd", x"03", x"fe", x"ff", x"ff", x"fd", x"00",
    x"fc", x"00", x"fd", x"fa", x"04", x"fc", x"04", x"fa",
    x"fd", x"fc", x"fa", x"ff", x"04", x"f8", x"00", x"fd",
    x"01", x"02", x"00", x"fa", x"fd", x"fc", x"02", x"fc",
    x"fe", x"00", x"fe", x"fb", x"03", x"fd", x"fc", x"fd",
    x"f9", x"02", x"02", x"01", x"01", x"03", x"00", x"01",
    x"fc", x"01", x"fc", x"04", x"fa", x"01", x"fa", x"04",
    x"2e", x"15", x"05", x"35", x"2c", x"f7", x"3f", x"20",
    x"01", x"16", x"db", x"07", x"06", x"fe", x"10", x"1a",
    x"e3", x"ec", x"16", x"f2", x"f9", x"f3", x"c0", x"e8",
    x"eb", x"ef", x"08", x"0a", x"16", x"35", x"30", x"12",
    x"22", x"33", x"16", x"3c", x"f9", x"da", x"01", x"22",
    x"06", x"10", x"07", x"10", x"32", x"c6", x"e3", x"af",
    x"13", x"bb", x"e1", x"00", x"ac", x"a5", x"06", x"0a",
    x"01", x"f5", x"0c", x"00", x"d8", x"0e", x"07", x"ec",
    x"06", x"65", x"ee", x"fc", x"42", x"fe", x"21", x"08",
    x"e9", x"fd", x"ea", x"e2", x"f4", x"17", x"07", x"03",
    x"fd", x"15", x"26", x"f6", x"93", x"cd", x"ee", x"7d",
    x"e6", x"da", x"2d", x"23", x"3c", x"78", x"ff", x"20",
    x"44", x"b5", x"22", x"00", x"01", x"1e", x"11", x"e8",
    x"f0", x"0d", x"bd", x"d4", x"04", x"ef", x"ec", x"18",
    x"ef", x"cf", x"25", x"c3", x"bb", x"b9", x"cf", x"84",
    x"b5", x"95", x"8c", x"a6", x"b5", x"df", x"42", x"35",
    x"11", x"f7", x"e2", x"e5", x"26", x"e8", x"2d", x"10",
    x"fd", x"f5", x"1a", x"0c", x"28", x"3f", x"27", x"08",
    x"af", x"fe", x"e4", x"a6", x"ea", x"ce", x"c0", x"a5",
    x"32", x"fb", x"04", x"fb", x"fc", x"05", x"fb", x"02",
    x"01", x"ff", x"e7", x"03", x"f6", x"ae", x"b0", x"c6",
    x"fb", x"ea", x"0a", x"b3", x"b8", x"cf", x"e3", x"c9",
    x"b2", x"8b", x"f1", x"ec", x"0a", x"05", x"10", x"31",
    x"09", x"03", x"2a", x"01", x"0f", x"18", x"24", x"f2",
    x"16", x"da", x"b7", x"b4", x"d6", x"01", x"20", x"0f",
    x"da", x"ee", x"fa", x"f5", x"be", x"e3", x"eb", x"8e",
    x"e4", x"bb", x"f0", x"fe", x"da", x"dd", x"f9", x"15",
    x"ad", x"ea", x"f2", x"17", x"f9", x"0e", x"ad", x"d7",
    x"0e", x"3c", x"2e", x"1b", x"4f", x"27", x"2d", x"4b",
    x"17", x"08", x"ea", x"fc", x"ff", x"cf", x"cd", x"a1",
    x"09", x"cb", x"e8", x"00", x"fa", x"02", x"06", x"fe",
    x"01", x"ff", x"fc", x"f8", x"f0", x"11", x"21", x"fa",
    x"07", x"fe", x"fd", x"0c", x"0c", x"02", x"0b", x"68",
    x"02", x"0d", x"3f", x"2f", x"5f", x"11", x"ff", x"e6",
    x"01", x"f2", x"b6", x"ec", x"ff", x"04", x"1b", x"24",
    x"02", x"12", x"0b", x"ff", x"fc", x"f4", x"d8", x"aa",
    x"0a", x"1d", x"2f", x"1f", x"07", x"26", x"57", x"25",
    x"16", x"e9", x"0d", x"e8", x"d9", x"da", x"ae", x"da",
    x"c8", x"b3", x"34", x"43", x"67", x"4e", x"2e", x"15",
    x"37", x"f3", x"fc", x"de", x"0b", x"fd", x"09", x"09",
    x"f2", x"0f", x"f3", x"f8", x"f7", x"03", x"02", x"f6",
    x"fa", x"fd", x"06", x"04", x"fb", x"f3", x"21", x"2d",
    x"10", x"0a", x"07", x"06", x"18", x"23", x"26", x"c6",
    x"e9", x"f0", x"a9", x"f5", x"79", x"bd", x"16", x"1d",
    x"02", x"0a", x"0d", x"02", x"f3", x"1c", x"ee", x"29",
    x"04", x"00", x"02", x"ff", x"02", x"03", x"04", x"02",
    x"00", x"f1", x"d6", x"fd", x"02", x"d5", x"dc", x"10",
    x"d6", x"ea", x"05", x"d1", x"f6", x"ed", x"ba", x"b8",
    x"06", x"89", x"6d", x"d8", x"e0", x"ed", x"ed", x"ed",
    x"e0", x"0e", x"c6", x"00", x"cb", x"e1", x"d8", x"ea",
    x"cb", x"dd", x"db", x"b0", x"b3", x"30", x"36", x"30",
    x"f0", x"11", x"e2", x"da", x"c5", x"ec", x"e4", x"17",
    x"cf", x"aa", x"fa", x"72", x"b6", x"fb", x"db", x"fc",
    x"e2", x"c1", x"b6", x"a0", x"98", x"0e", x"15", x"d4",
    x"fc", x"fd", x"fc", x"01", x"fe", x"05", x"fe", x"fe",
    x"02", x"fd", x"04", x"03", x"00", x"02", x"06", x"fd",
    x"fd", x"fe", x"38", x"2c", x"1a", x"1c", x"3f", x"18",
    x"e2", x"35", x"11", x"f4", x"f9", x"e0", x"1a", x"d5",
    x"cc", x"0d", x"f8", x"33", x"d7", x"ed", x"7d", x"c2",
    x"a5", x"9e", x"01", x"25", x"d1", x"cf", x"f8", x"f9",
    x"c9", x"09", x"2b", x"b5", x"00", x"f5", x"14", x"1d",
    x"18", x"cd", x"f9", x"ec", x"b6", x"ea", x"1b", x"b0",
    x"ef", x"ff", x"38", x"f7", x"0d", x"4b", x"e4", x"e5",
    x"2a", x"1b", x"f7", x"02", x"f8", x"cc", x"b4", x"f8",
    x"e4", x"5d", x"44", x"10", x"4c", x"3c", x"00", x"1e",
    x"29", x"1b", x"0b", x"eb", x"b1", x"2a", x"41", x"44",
    x"42", x"3e", x"38", x"1c", x"fa", x"22", x"ff", x"0e",
    x"02", x"55", x"08", x"fb", x"02", x"04", x"d7", x"0e",
    x"01", x"f3", x"0b", x"dd", x"f3", x"d5", x"e1", x"f1",
    x"09", x"12", x"bd", x"ec", x"e8", x"ca", x"08", x"1d",
    x"35", x"03", x"02", x"16", x"67", x"de", x"24", x"26",
    x"26", x"24", x"0e", x"e9", x"19", x"1f", x"e5", x"de",
    x"e6", x"03", x"7d", x"d8", x"f3", x"dd", x"bf", x"aa",
    x"b2", x"fc", x"f2", x"03", x"7c", x"f3", x"c1", x"ef",
    x"f3", x"a1", x"ad", x"cf", x"05", x"a6", x"af", x"db",
    x"d1", x"2f", x"c6", x"e4", x"d5", x"00", x"ad", x"ec",
    x"05", x"1b", x"05", x"0c", x"f0", x"10", x"22", x"98",
    x"af", x"9d", x"0b", x"3d", x"25", x"ea", x"fa", x"09",
    x"2c", x"ec", x"a9", x"52", x"56", x"f8", x"16", x"31",
    x"23", x"29", x"02", x"fe", x"f6", x"0e", x"15", x"08",
    x"fc", x"41", x"26", x"23", x"31", x"d1", x"e2", x"0a",
    x"dd", x"ec", x"24", x"11", x"0b", x"51", x"aa", x"c0",
    x"ce", x"bb", x"a4", x"f2", x"ff", x"1a", x"5a", x"cc",
    x"fa", x"46", x"0a", x"f9", x"0e", x"d3", x"c0", x"fe",
    x"f9", x"10", x"1e", x"5b", x"19", x"02", x"3d", x"04",
    x"f3", x"12", x"db", x"20", x"0e", x"ec", x"da", x"00",
    x"a8", x"ce", x"dc", x"c8", x"ca", x"f6", x"17", x"3e",
    x"fe", x"15", x"28", x"f4", x"f2", x"0a", x"ed", x"d7",
    x"ee", x"1f", x"32", x"13", x"2a", x"24", x"1d", x"98",
    x"ee", x"18", x"04", x"08", x"0f", x"f1", x"f0", x"fe",
    x"24", x"43", x"32", x"ef", x"c7", x"90", x"d7", x"d7",
    x"d0", x"fc", x"fd", x"05", x"02", x"00", x"05", x"03",
    x"03", x"01", x"35", x"1c", x"27", x"f5", x"21", x"0f",
    x"24", x"1d", x"f7", x"ee", x"e0", x"f1", x"e2", x"f9",
    x"2e", x"f5", x"fe", x"e1", x"e9", x"fb", x"fa", x"21",
    x"29", x"2a", x"3e", x"14", x"2b", x"f9", x"de", x"f4",
    x"8b", x"9c", x"f4", x"b3", x"dc", x"c9", x"06", x"0c",
    x"03", x"c9", x"96", x"95", x"7a", x"a4", x"8e", x"0c",
    x"ee", x"fc", x"dd", x"cf", x"c6", x"0b", x"f7", x"f9",
    x"0a", x"59", x"11", x"46", x"b2", x"ed", x"22", x"05",
    x"b7", x"04", x"fb", x"42", x"2e", x"1b", x"19", x"05",
    x"f4", x"d4", x"e5", x"f9", x"f5", x"ab", x"aa", x"8e",
    x"ae", x"14", x"f8", x"06", x"05", x"fb", x"01", x"03",
    x"fc", x"0b", x"05", x"07", x"e0", x"f7", x"08", x"f9",
    x"27", x"16", x"e7", x"19", x"03", x"08", x"05", x"07",
    x"aa", x"04", x"20", x"35", x"47", x"28", x"16", x"1c",
    x"09", x"32", x"2a", x"0d", x"23", x"1c", x"31", x"f8",
    x"fc", x"09", x"21", x"2c", x"2e", x"e0", x"1d", x"2f",
    x"11", x"14", x"1c", x"0a", x"0a", x"0e", x"e7", x"0b",
    x"fd", x"fb", x"d7", x"0a", x"f3", x"39", x"d0", x"05",
    x"2e", x"39", x"3e", x"29", x"2d", x"60", x"29", x"fd",
    x"7f", x"dd", x"e2", x"de", x"01", x"25", x"18", x"42",
    x"1b", x"ac", x"ee", x"04", x"0a", x"04", x"06", x"0c",
    x"08", x"fb", x"10", x"05", x"05", x"ff", x"28", x"29",
    x"f8", x"18", x"ed", x"f0", x"06", x"36", x"e6", x"ca",
    x"01", x"f9", x"16", x"31", x"d3", x"10", x"fe", x"f0",
    x"f9", x"1f", x"cf", x"f7", x"f7", x"ef", x"08", x"0c",
    x"07", x"fb", x"fc", x"fd", x"02", x"05", x"02", x"05",
    x"00", x"3d", x"04", x"02", x"fc", x"0f", x"23", x"ca",
    x"0f", x"f5", x"53", x"fd", x"09", x"ec", x"12", x"2e",
    x"db", x"e7", x"df", x"ef", x"19", x"2f", x"ea", x"23",
    x"0c", x"1e", x"aa", x"a3", x"ca", x"e6", x"e6", x"ef",
    x"d5", x"b8", x"29", x"18", x"0a", x"fd", x"12", x"ff",
    x"2c", x"10", x"33", x"70", x"89", x"78", x"42", x"1b",
    x"27", x"e2", x"0a", x"0e", x"08", x"0c", x"1b", x"e4",
    x"df", x"ee", x"c0", x"e7", x"d9", x"fd", x"f2", x"d6",
    x"01", x"08", x"01", x"f7", x"fe", x"02", x"fe", x"02",
    x"fd", x"fd", x"08", x"fb", x"07", x"04", x"01", x"09",
    x"fc", x"fa", x"ea", x"e0", x"d8", x"86", x"91", x"ca",
    x"c2", x"ec", x"f1", x"0c", x"2b", x"01", x"1a", x"f9",
    x"10", x"02", x"f1", x"0f", x"e6", x"df", x"f9", x"08",
    x"e7", x"fb", x"1f", x"27", x"50", x"22", x"0e", x"fd",
    x"fc", x"ec", x"f6", x"aa", x"c8", x"29", x"09", x"db",
    x"11", x"e9", x"e1", x"c3", x"25", x"0f", x"10", x"3c",
    x"35", x"18", x"20", x"13", x"1c", x"18", x"35", x"1f",
    x"24", x"39", x"f9", x"1a", x"f3", x"33", x"ea", x"07",
    x"06", x"2e", x"18", x"15", x"f7", x"38", x"0a", x"3a",
    x"2b", x"26", x"f0", x"d5", x"e7", x"35", x"11", x"43",
    x"dd", x"1a", x"1f", x"21", x"fc", x"df", x"0f", x"c4",
    x"c2", x"c7", x"d8", x"cd", x"26", x"31", x"2b", x"15",
    x"12", x"1e", x"e9", x"00", x"02", x"1c", x"13", x"06",
    x"12", x"04", x"13", x"c8", x"13", x"46", x"25", x"3a",
    x"ff", x"16", x"d7", x"0a", x"04", x"d9", x"00", x"22",
    x"08", x"3d", x"19", x"1c", x"01", x"18", x"f2", x"1b",
    x"fd", x"e7", x"dc", x"e9", x"f6", x"17", x"d5", x"f2",
    x"2b", x"00", x"33", x"40", x"a8", x"f6", x"2f", x"ff",
    x"e0", x"f5", x"b2", x"e2", x"e0", x"21", x"14", x"e3",
    x"01", x"1b", x"0c", x"d5", x"c2", x"a7", x"2c", x"14",
    x"a4", x"20", x"37", x"05", x"fa", x"fc", x"0a", x"d4",
    x"fd", x"12", x"0e", x"3b", x"4c", x"cc", x"0a", x"2e",
    x"a7", x"d1", x"da", x"7d", x"a8", x"b8", x"31", x"0e",
    x"16", x"95", x"e0", x"e5", x"f7", x"09", x"0e", x"9b",
    x"55", x"20", x"23", x"ff", x"dd", x"00", x"da", x"ef",
    x"38", x"14", x"28", x"1c", x"16", x"43", x"34", x"2a",
    x"31", x"de", x"b3", x"dd", x"f7", x"ff", x"e1", x"18",
    x"e6", x"0a", x"b7", x"7b", x"94", x"08", x"9a", x"d2",
    x"fb", x"11", x"0a", x"3c", x"22", x"f9", x"40", x"cb",
    x"d5", x"e6", x"be", x"c2", x"2b", x"36", x"0b", x"d7",
    x"ee", x"08", x"33", x"28", x"ee", x"f2", x"e8", x"a7",
    x"08", x"f9", x"e1", x"1e", x"14", x"d6", x"0e", x"fe",
    x"2c", x"66", x"5c", x"16", x"35", x"24", x"ec", x"ea",
    x"1c", x"0d", x"23", x"fc", x"b2", x"4a", x"10", x"d2",
    x"1b", x"2b", x"3e", x"06", x"20", x"3e", x"22", x"1c",
    x"1d", x"fd", x"fd", x"fe", x"04", x"fe", x"fb", x"02",
    x"ff", x"03", x"04", x"9b", x"c1", x"0e", x"25", x"0a",
    x"f7", x"f1", x"f8", x"f9", x"f2", x"16", x"c2", x"18",
    x"06", x"1b", x"36", x"cf", x"0f", x"f7", x"df", x"22",
    x"f9", x"f2", x"e4", x"ef", x"cb", x"a4", x"f1", x"f4",
    x"bc", x"e5", x"fc", x"f5", x"c3", x"b7", x"fa", x"e8",
    x"da", x"eb", x"ee", x"f5", x"d9", x"fe", x"eb", x"fe",
    x"1d", x"ff", x"e2", x"3a", x"2d", x"e5", x"0f", x"13",
    x"35", x"17", x"06", x"0e", x"26", x"39", x"91", x"29",
    x"2f", x"d9", x"f0", x"cf", x"06", x"fd", x"01", x"b1",
    x"e5", x"fe", x"ae", x"ea", x"1c", x"b1", x"09", x"1d",
    x"6c", x"7d", x"5d", x"f8", x"01", x"05", x"01", x"03",
    x"ff", x"00", x"ff", x"04", x"fc", x"12", x"1c", x"ef",
    x"29", x"1d", x"09", x"fa", x"30", x"14", x"0c", x"fd",
    x"f2", x"c8", x"b6", x"06", x"9d", x"ff", x"e7", x"dc",
    x"e0", x"32", x"11", x"fd", x"3a", x"ea", x"df", x"1a",
    x"4b", x"58", x"22", x"14", x"36", x"c4", x"e8", x"04",
    x"1c", x"29", x"fa", x"f4", x"fc", x"2b", x"f5", x"f8",
    x"fb", x"ec", x"ef", x"07", x"f9", x"fb", x"06", x"01",
    x"f5", x"03", x"23", x"33", x"0c", x"1b", x"fa", x"fb",
    x"ef", x"e4", x"b0", x"e6", x"e9", x"23", x"ec", x"f0",
    x"15", x"7a", x"14", x"14", x"00", x"f6", x"01", x"f9",
    x"00", x"fd", x"03", x"fd", x"fc", x"f2", x"dd", x"bc",
    x"1f", x"e1", x"e7", x"2e", x"f1", x"c1", x"e5", x"dc",
    x"ef", x"48", x"18", x"0b", x"fc", x"12", x"25", x"04",
    x"08", x"e4", x"e9", x"fb", x"e0", x"c2", x"20", x"04",
    x"fe", x"fe", x"fc", x"02", x"04", x"fb", x"02", x"fc",
    x"fc", x"cf", x"c5", x"ed", x"25", x"cb", x"ea", x"46",
    x"ee", x"01", x"14", x"f7", x"f4", x"ce", x"ec", x"15",
    x"c4", x"db", x"3e", x"0e", x"03", x"f7", x"69", x"55",
    x"2d", x"47", x"fc", x"15", x"ed", x"14", x"ca", x"35",
    x"fd", x"00", x"f9", x"26", x"0b", x"0d", x"03", x"19",
    x"f3", x"06", x"32", x"ef", x"12", x"42", x"06", x"bd",
    x"32", x"d6", x"c8", x"00", x"fd", x"f3", x"f2", x"ee",
    x"d9", x"f9", x"09", x"0c", x"01", x"fc", x"17", x"0d",
    x"06", x"fc", x"03", x"fb", x"ff", x"fe", x"08", x"05",
    x"06", x"fa", x"ff", x"ff", x"fb", x"fd", x"01", x"fc",
    x"fc", x"fa", x"d7", x"04", x"04", x"11", x"37", x"3d",
    x"38", x"3c", x"40", x"dc", x"21", x"37", x"f1", x"f7",
    x"3e", x"09", x"ec", x"94", x"a1", x"da", x"f8", x"cc",
    x"cf", x"f1", x"dd", x"f5", x"c9", x"2e", x"25", x"3e",
    x"d2", x"32", x"2a", x"be", x"87", x"c1", x"bf", x"fa",
    x"f4", x"0c", x"00", x"0c", x"c7", x"cb", x"de", x"42",
    x"43", x"11", x"f0", x"da", x"ec", x"0f", x"ca", x"d8",
    x"09", x"ea", x"dd", x"da", x"b2", x"c1", x"f4", x"06",
    x"fe", x"e7", x"20", x"3c", x"d3", x"ec", x"14", x"e0",
    x"a1", x"fc", x"f9", x"ed", x"00", x"fb", x"b1", x"bc",
    x"37", x"f4", x"ab", x"00", x"f4", x"01", x"1a", x"f2",
    x"dd", x"bf", x"d3", x"8f", x"24", x"41", x"28", x"e6",
    x"d8", x"f1", x"09", x"0c", x"eb", x"ff", x"34", x"26",
    x"e1", x"e7", x"fa", x"d1", x"a9", x"df", x"6f", x"de",
    x"e4", x"cb", x"d5", x"07", x"cb", x"09", x"03", x"11",
    x"24", x"17", x"d8", x"f4", x"3d", x"d5", x"e5", x"d5",
    x"d3", x"0d", x"fd", x"f5", x"30", x"bd", x"1f", x"4c",
    x"1c", x"d2", x"fe", x"11", x"d3", x"f4", x"34", x"f0",
    x"33", x"14", x"76", x"29", x"71", x"a5", x"ed", x"a4",
    x"9a", x"b6", x"8d", x"2e", x"1f", x"01", x"09", x"e4",
    x"09", x"ff", x"f2", x"38", x"e2", x"37", x"0f", x"00",
    x"f2", x"07", x"fb", x"f2", x"18", x"fc", x"e7", x"19",
    x"d9", x"03", x"5f", x"14", x"17", x"0a", x"0a", x"fd",
    x"11", x"0a", x"13", x"13", x"1f", x"25", x"38", x"d2",
    x"0a", x"0b", x"b4", x"cf", x"cd", x"f8", x"14", x"19",
    x"cd", x"fa", x"fc", x"f6", x"f0", x"b7", x"11", x"04",
    x"f4", x"e8", x"f1", x"12", x"c4", x"e0", x"05", x"1c",
    x"23", x"38", x"45", x"12", x"26", x"07", x"01", x"ff",
    x"02", x"c7", x"cc", x"10", x"06", x"1a", x"25", x"d5",
    x"d1", x"44", x"d5", x"d3", x"f4", x"06", x"e2", x"0b",
    x"06", x"2a", x"fa", x"16", x"05", x"c4", x"e6", x"24",
    x"f0", x"cf", x"f5", x"f0", x"01", x"01", x"28", x"37",
    x"ea", x"be", x"c8", x"f0", x"b0", x"95", x"d5", x"bb",
    x"c7", x"bb", x"a0", x"a0", x"96", x"b9", x"b6", x"07",
    x"19", x"e2", x"e9", x"21", x"0e", x"2a", x"18", x"25",
    x"12", x"ff", x"05", x"fd", x"03", x"02", x"fd", x"02",
    x"ff", x"ff", x"28", x"0c", x"49", x"2a", x"1a", x"3c",
    x"d2", x"e4", x"b2", x"e6", x"25", x"20", x"e9", x"12",
    x"2c", x"2b", x"fe", x"18", x"e0", x"f1", x"06", x"e7",
    x"f5", x"09", x"23", x"0c", x"f5", x"fd", x"0b", x"fa",
    x"ea", x"f7", x"e2", x"e0", x"f9", x"09", x"3f", x"2e",
    x"f3", x"21", x"19", x"1c", x"ee", x"eb", x"cf", x"bc",
    x"d6", x"ff", x"ed", x"06", x"d6", x"18", x"ec", x"fe",
    x"f4", x"2a", x"fb", x"0c", x"27", x"e2", x"13", x"06",
    x"cc", x"fa", x"eb", x"0c", x"cb", x"e5", x"00", x"28",
    x"07", x"1a", x"2c", x"ed", x"c7", x"08", x"0b", x"04",
    x"07", x"12", x"1d", x"fb", x"fb", x"fe", x"ff", x"fc",
    x"fb", x"fb", x"fe", x"02", x"00", x"3b", x"22", x"f8",
    x"f6", x"d4", x"fb", x"e4", x"dd", x"dd", x"03", x"17",
    x"f5", x"d1", x"cb", x"0f", x"1d", x"c6", x"bf", x"d1",
    x"f5", x"dd", x"f0", x"0d", x"e5", x"f6", x"20", x"fe",
    x"db", x"10", x"d5", x"af", x"be", x"f4", x"eb", x"0b",
    x"ce", x"f9", x"ff", x"fd", x"2b", x"d0", x"25", x"3e",
    x"c1", x"ed", x"fa", x"e6", x"f3", x"c3", x"ef", x"e4",
    x"cf", x"01", x"ce", x"bc", x"0e", x"16", x"0d", x"07",
    x"ec", x"19", x"df", x"d4", x"25", x"12", x"01", x"cc",
    x"82", x"3f", x"21", x"2d", x"f9", x"fb", x"fc", x"00",
    x"fd", x"03", x"fe", x"f7", x"01", x"eb", x"f4", x"ea",
    x"c2", x"0d", x"1b", x"c2", x"1d", x"30", x"1d", x"e4",
    x"e2", x"16", x"a7", x"b8", x"4d", x"b1", x"87", x"32",
    x"e7", x"ff", x"2a", x"03", x"b9", x"38", x"f9", x"0f",
    x"fd", x"03", x"fe", x"fd", x"01", x"03", x"05", x"06",
    x"01", x"e8", x"a0", x"b3", x"f7", x"a9", x"61", x"eb",
    x"f9", x"01", x"0d", x"1c", x"f8", x"18", x"f9", x"c3",
    x"08", x"2d", x"f5", x"31", x"d9", x"0d", x"12", x"5e",
    x"c9", x"20", x"10", x"23", x"cc", x"cf", x"cd", x"02",
    x"ef", x"18", x"e1", x"0d", x"36", x"1d", x"b9", x"ea",
    x"3b", x"29", x"1a", x"04", x"07", x"17", x"2c", x"6b",
    x"36", x"4a", x"51", x"0f", x"fb", x"ed", x"e8", x"f2",
    x"e8", x"1e", x"02", x"1b", x"3d", x"11", x"1d", x"23",
    x"fc", x"fd", x"01", x"03", x"04", x"fc", x"fe", x"04",
    x"05", x"fd", x"01", x"fd", x"ff", x"fc", x"02", x"05",
    x"02", x"02", x"48", x"64", x"2e", x"29", x"f5", x"26",
    x"13", x"04", x"09", x"21", x"0e", x"ad", x"2d", x"2a",
    x"21", x"39", x"09", x"97", x"cd", x"ee", x"0c", x"14",
    x"c7", x"0d", x"e1", x"ab", x"f5", x"ce", x"c1", x"d2",
    x"eb", x"eb", x"ef", x"f2", x"f9", x"07", x"fa", x"0d",
    x"31", x"76", x"16", x"e7", x"18", x"d6", x"a7", x"c5",
    x"bb", x"e7", x"ed", x"d9", x"ea", x"35", x"f1", x"10",
    x"1b", x"16", x"17", x"0f", x"0d", x"bd", x"08", x"fc",
    x"93", x"02", x"fc", x"ca", x"1e", x"2c", x"09", x"f1",
    x"16", x"4f", x"e9", x"f9", x"db", x"dd", x"12", x"fe",
    x"e2", x"ec", x"09", x"f5", x"da", x"dd", x"2a", x"20",
    x"08", x"0f", x"f3", x"c7", x"df", x"fa", x"e2", x"09",
    x"d8", x"ee", x"29", x"12", x"13", x"06", x"f2", x"16",
    x"01", x"09", x"3b", x"ef", x"35", x"48", x"03", x"eb",
    x"fd", x"17", x"2b", x"fc", x"12", x"0a", x"fd", x"e2",
    x"af", x"18", x"0c", x"27", x"53", x"18", x"1a", x"11",
    x"0e", x"31", x"18", x"1b", x"17", x"f8", x"43", x"26",
    x"3e", x"28", x"f3", x"eb", x"b8", x"fe", x"08", x"f4",
    x"f7", x"e4", x"fb", x"10", x"2f", x"e5", x"0e", x"39",
    x"0b", x"f6", x"11", x"0c", x"0b", x"19", x"30", x"38",
    x"0a", x"f8", x"f3", x"ea", x"d8", x"f4", x"e1", x"aa",
    x"cb", x"e1", x"d2", x"a7", x"ee", x"fe", x"12", x"30",
    x"b2", x"17", x"30", x"dc", x"f1", x"ee", x"cd", x"0d",
    x"2c", x"43", x"22", x"06", x"1d", x"09", x"20", x"fa",
    x"05", x"13", x"32", x"09", x"12", x"25", x"2f", x"2c",
    x"11", x"fa", x"1d", x"e9", x"0e", x"ea", x"28", x"14",
    x"f1", x"d9", x"be", x"e4", x"97", x"a3", x"f6", x"9a",
    x"aa", x"dc", x"44", x"2f", x"39", x"47", x"28", x"47",
    x"08", x"3d", x"32", x"08", x"05", x"f7", x"f3", x"03",
    x"0b", x"2c", x"11", x"18", x"ef", x"a0", x"d4", x"3e",
    x"a8", x"b6", x"2b", x"b0", x"87", x"c9", x"e7", x"19",
    x"ce", x"ef", x"e7", x"b3", x"e5", x"a2", x"ee", x"87",
    x"b2", x"7a", x"46", x"79", x"d0", x"93", x"96", x"50",
    x"2a", x"29", x"27", x"1b", x"14", x"16", x"0c", x"0d",
    x"c3", x"d4", x"e4", x"65", x"f4", x"20", x"13", x"0d",
    x"4f", x"02", x"fb", x"00", x"fd", x"fd", x"04", x"05",
    x"fc", x"03", x"cf", x"ba", x"db", x"9a", x"60", x"78",
    x"fc", x"e5", x"e0", x"e3", x"01", x"e8", x"d3", x"25",
    x"0f", x"ab", x"03", x"1c", x"20", x"26", x"31", x"f1",
    x"0b", x"fe", x"d0", x"11", x"39", x"ed", x"9a", x"fd",
    x"95", x"ad", x"f3", x"0e", x"f8", x"c9", x"e9", x"f1",
    x"0e", x"eb", x"fe", x"fa", x"3d", x"2d", x"2d", x"a7",
    x"be", x"e7", x"36", x"ff", x"30", x"20", x"d9", x"0c",
    x"2b", x"21", x"15", x"0b", x"14", x"eb", x"3f", x"2d",
    x"08", x"28", x"43", x"17", x"02", x"16", x"0b", x"cb",
    x"1c", x"31", x"cf", x"fb", x"f8", x"dc", x"db", x"f9",
    x"d9", x"d0", x"ae", x"03", x"ff", x"fe", x"04", x"fb",
    x"f8", x"05", x"01", x"ff", x"c6", x"e5", x"c4", x"d3",
    x"9b", x"ae", x"d0", x"c2", x"b3", x"f7", x"02", x"3b",
    x"1f", x"1e", x"31", x"2f", x"08", x"28", x"0c", x"e7",
    x"fa", x"bd", x"cb", x"d3", x"d3", x"d7", x"fa", x"eb",
    x"b4", x"d7", x"b9", x"ad", x"cd", x"db", x"af", x"6d",
    x"30", x"1f", x"12", x"14", x"05", x"fd", x"14", x"05",
    x"0a", x"c3", x"04", x"3b", x"86", x"91", x"c4", x"ee",
    x"e8", x"e4", x"4f", x"42", x"49", x"30", x"26", x"20",
    x"0e", x"0d", x"20", x"36", x"36", x"30", x"19", x"b9",
    x"d4", x"43", x"d1", x"ce", x"10", x"05", x"04", x"0a",
    x"01", x"10", x"0c", x"05", x"06", x"62", x"3b", x"f9",
    x"60", x"0d", x"ff", x"2e", x"f4", x"07", x"15", x"16",
    x"19", x"3e", x"fd", x"0a", x"3e", x"ff", x"07", x"fe",
    x"1a", x"03", x"1f", x"1a", x"15", x"27", x"15", x"0f",
    x"00", x"fc", x"fb", x"fd", x"ff", x"01", x"02", x"01",
    x"fe", x"01", x"dc", x"db", x"d7", x"ee", x"f4", x"ec",
    x"03", x"df", x"2f", x"fb", x"dd", x"39", x"f9", x"00",
    x"4c", x"fc", x"d2", x"3c", x"e4", x"e9", x"bc", x"d4",
    x"eb", x"10", x"cb", x"e3", x"26", x"3f", x"0b", x"05",
    x"f5", x"e2", x"d9", x"eb", x"10", x"da", x"07", x"1e",
    x"0a", x"11", x"0b", x"d1", x"e9", x"fa", x"be", x"e7",
    x"14", x"ce", x"c6", x"f2", x"f4", x"18", x"04", x"be",
    x"b9", x"2d", x"c3", x"8a", x"fb", x"ee", x"df", x"fd",
    x"04", x"05", x"05", x"fc", x"04", x"fd", x"03", x"fe",
    x"fc", x"03", x"fa", x"ff", x"00", x"00", x"fe", x"02",
    x"fc", x"06", x"07", x"e0", x"f6", x"1b", x"f7", x"0a",
    x"0e", x"2a", x"10", x"ff", x"f4", x"e2", x"10", x"f4",
    x"c3", x"db", x"fa", x"c3", x"ea", x"d5", x"cf", x"ab",
    x"b6", x"af", x"a6", x"ee", x"15", x"9f", x"b5", x"bc",
    x"bf", x"b9", x"c9", x"2e", x"ce", x"d3", x"bb", x"e2",
    x"f6", x"9e", x"f1", x"e0", x"e9", x"02", x"03", x"db",
    x"22", x"0c", x"23", x"fc", x"fc", x"38", x"0f", x"f6",
    x"13", x"1b", x"1d", x"f3", x"ef", x"e8", x"0d", x"14",
    x"15", x"d5", x"ca", x"ef", x"a5", x"e2", x"f1", x"b8",
    x"e7", x"e9", x"68", x"16", x"ed", x"51", x"20", x"16",
    x"25", x"37", x"2c", x"d6", x"7c", x"a6", x"ff", x"c8",
    x"b6", x"f1", x"e0", x"dd", x"fa", x"11", x"f2", x"14",
    x"f6", x"c9", x"e3", x"19", x"e6", x"05", x"04", x"0e",
    x"02", x"18", x"cb", x"42", x"30", x"c5", x"1d", x"f0",
    x"13", x"2a", x"31", x"4b", x"06", x"15", x"0d", x"ec",
    x"2c", x"55", x"39", x"38", x"32", x"fd", x"2b", x"07",
    x"fc", x"f7", x"00", x"f7", x"fd", x"03", x"00", x"fd",
    x"01", x"fc", x"f6", x"04", x"02", x"f7", x"fc", x"f8",
    x"03", x"fb", x"fb", x"fd", x"ff", x"02", x"ff", x"ff",
    x"01", x"01", x"f9", x"fa", x"f9", x"fb", x"fd", x"fb",
    x"fa", x"f8", x"fb", x"f9", x"ff", x"01", x"fb", x"00",
    x"f7", x"f9", x"fb", x"00", x"f9", x"fa", x"fb", x"ff",
    x"fb", x"f8", x"fb", x"fc", x"01", x"02", x"fd", x"f8",
    x"fc", x"ff", x"fd", x"f6", x"ff", x"fc", x"fd", x"fb",
    x"03", x"00", x"fc", x"fa", x"fc", x"f8", x"00", x"f7",
    x"fd", x"fb", x"ff", x"ff", x"01", x"ff", x"fe", x"fe",
    x"02", x"01", x"f4", x"03", x"02", x"00", x"ff", x"fb",
    x"01", x"02", x"fa", x"fd", x"f7", x"fd", x"00", x"02",
    x"01", x"fc", x"fc", x"01", x"fd", x"f8", x"fc", x"f7",
    x"fb", x"fd", x"fa", x"01", x"02", x"fd", x"fd", x"fd",
    x"fc", x"01", x"03", x"fe", x"f7", x"fb", x"00", x"fd",
    x"fc", x"fb", x"f8", x"fb", x"ff", x"fb", x"fb", x"ff",
    x"fa", x"fa", x"ff", x"fd", x"fd", x"f7", x"f8", x"fb",
    x"f7", x"f8", x"f8", x"fb", x"f8", x"01", x"00", x"00",
    x"fe", x"f9", x"02", x"f8", x"00", x"07", x"01", x"fb",
    x"01", x"00", x"ff", x"fb", x"05", x"04", x"01", x"01",
    x"02", x"00", x"f9", x"fb", x"ff", x"fb", x"fe", x"fc",
    x"01", x"01", x"f7", x"00", x"ff", x"04", x"01", x"fd",
    x"03", x"fb", x"02", x"02", x"fc", x"fd", x"fe", x"fe",
    x"fb", x"fa", x"01", x"fb", x"fe", x"fb", x"02", x"ff",
    x"fd", x"f8", x"ff", x"fb", x"01", x"fe", x"fd", x"fd",
    x"fb", x"fe", x"f8", x"00", x"f8", x"f8", x"fe", x"ff",
    x"f9", x"fc", x"fe", x"fe", x"fe", x"fd", x"04", x"fc",
    x"fc", x"fb", x"ff", x"03", x"fe", x"01", x"fc", x"04",
    x"01", x"fc", x"00", x"fe", x"04", x"00", x"f8", x"ff",
    x"fc", x"fc", x"fb", x"fa", x"f9", x"04", x"00", x"fb",
    x"fc", x"fe", x"00", x"fd", x"fd", x"00", x"02", x"01",
    x"00", x"01", x"04", x"00", x"00", x"ff", x"fc", x"00",
    x"f7", x"f8", x"ff", x"fa", x"f9", x"f8", x"fd", x"00",
    x"01", x"f6", x"fa", x"ff", x"ff", x"fe", x"fc", x"f7",
    x"00", x"fc", x"ff", x"fb", x"01", x"f6", x"00", x"02",
    x"04", x"01", x"fd", x"f8", x"02", x"fa", x"ff", x"fe",
    x"f9", x"02", x"fe", x"f9", x"fb", x"00", x"f7", x"f9",
    x"fc", x"01", x"f8", x"00", x"fd", x"f7", x"ff", x"fc",
    x"fe", x"00", x"ff", x"01", x"fa", x"03", x"ff", x"00",
    x"fa", x"fb", x"f7", x"fe", x"ff", x"00", x"f7", x"f6",
    x"ff", x"fc", x"fd", x"fa", x"ff", x"05", x"02", x"05",
    x"03", x"02", x"fb", x"01", x"fd", x"00", x"00", x"fc",
    x"fe", x"03", x"f7", x"00", x"fa", x"fe", x"04", x"ff",
    x"fc", x"ff", x"01", x"fb", x"00", x"01", x"f9", x"f8",
    x"fd", x"00", x"00", x"00", x"02", x"fb", x"00", x"f8",
    x"03", x"fe", x"03", x"05", x"04", x"fe", x"01", x"05",
    x"fe", x"fb", x"fc", x"fd", x"ff", x"03", x"00", x"00",
    x"fa", x"01", x"fc", x"00", x"fd", x"03", x"01", x"01",
    x"04", x"01", x"fa", x"fc", x"fb", x"fe", x"fc", x"fb",
    x"fd", x"fe", x"03", x"fe", x"fd", x"fd", x"02", x"fb",
    x"fe", x"ff", x"fc", x"02", x"00", x"00", x"00", x"01",
    x"fd", x"fd", x"fd", x"00", x"f8", x"fc", x"f6", x"f9",
    x"fb", x"fc", x"fe", x"ff", x"fe", x"00", x"f9", x"fc",
    x"f8", x"fc", x"fe", x"f7", x"fd", x"fe", x"f8", x"02",
    x"fd", x"05", x"00", x"fd", x"02", x"fd", x"fe", x"03",
    x"ff", x"02", x"00", x"02", x"02", x"fe", x"05", x"02",
    x"04", x"fc", x"fe", x"02", x"03", x"f7", x"ff", x"f7",
    x"01", x"00", x"03", x"fb", x"00", x"ff", x"f8", x"fb",
    x"fc", x"fc", x"fd", x"fd", x"fd", x"00", x"fe", x"f7",
    x"f4", x"f9", x"01", x"04", x"fd", x"fb", x"f4", x"00",
    x"fc", x"fd", x"01", x"f9", x"ff", x"ff", x"f7", x"f8",
    x"00", x"fd", x"fc", x"fe", x"f9", x"f7", x"01", x"01",
    x"fc", x"ff", x"04", x"fe", x"fd", x"fd", x"01", x"ff",
    x"04", x"fa", x"02", x"fc", x"f7", x"fb", x"f9", x"05",
    x"01", x"00", x"f6", x"f7", x"03", x"f8", x"fb", x"fc",
    x"f9", x"00", x"01", x"01", x"fb", x"01", x"00", x"00",
    x"01", x"f7", x"ff", x"ff", x"fb", x"03", x"fc", x"fb",
    x"00", x"fa", x"fa", x"fb", x"ff", x"ff", x"ff", x"00",
    x"00", x"06", x"fd", x"ff", x"fd", x"f9", x"fc", x"f6",
    x"00", x"ff", x"02", x"fd", x"f8", x"ff", x"fe", x"02",
    x"fb", x"00", x"02", x"02", x"01", x"04", x"fe", x"fe",
    x"fd", x"fc", x"fe", x"fb", x"fd", x"05", x"f9", x"ff",
    x"46", x"34", x"13", x"2b", x"35", x"fa", x"2d", x"17",
    x"03", x"f5", x"0a", x"0f", x"10", x"e6", x"f7", x"06",
    x"da", x"e0", x"ba", x"e4", x"f7", x"eb", x"db", x"cf",
    x"1c", x"d4", x"c2", x"fe", x"01", x"fd", x"17", x"4a",
    x"0d", x"08", x"f0", x"fc", x"dc", x"d8", x"ed", x"09",
    x"02", x"31", x"e3", x"1a", x"45", x"1d", x"23", x"46",
    x"19", x"d3", x"9b", x"0a", x"ec", x"b4", x"08", x"ea",
    x"f5", x"31", x"16", x"19", x"17", x"31", x"23", x"4f",
    x"0c", x"2a", x"b3", x"c3", x"f8", x"15", x"fb", x"0d",
    x"18", x"f8", x"00", x"00", x"e1", x"cd", x"fc", x"d9",
    x"14", x"23", x"12", x"2a", x"f2", x"bf", x"a3", x"b9",
    x"7a", x"ed", x"2d", x"16", x"2b", x"35", x"48", x"2b",
    x"0b", x"0c", x"27", x"24", x"d2", x"d7", x"bc", x"28",
    x"ff", x"02", x"32", x"0a", x"32", x"29", x"ba", x"1f",
    x"f7", x"d5", x"2b", x"db", x"9c", x"f8", x"c1", x"0e",
    x"de", x"ed", x"02", x"cc", x"ae", x"f5", x"29", x"14",
    x"02", x"d3", x"cb", x"d8", x"ea", x"c8", x"b6", x"1a",
    x"e2", x"0f", x"23", x"08", x"10", x"13", x"fb", x"fc",
    x"09", x"19", x"de", x"05", x"dc", x"da", x"cc", x"d6",
    x"ad", x"04", x"ff", x"fd", x"fe", x"05", x"fc", x"fd",
    x"00", x"01", x"10", x"00", x"13", x"f6", x"cf", x"ee",
    x"ea", x"d1", x"e8", x"05", x"f4", x"f8", x"16", x"e6",
    x"ea", x"c8", x"07", x"34", x"1b", x"f5", x"14", x"fa",
    x"fb", x"1d", x"17", x"ce", x"1e", x"39", x"1a", x"1e",
    x"16", x"19", x"23", x"e6", x"a6", x"fa", x"2a", x"36",
    x"34", x"0d", x"02", x"0b", x"07", x"08", x"ee", x"f6",
    x"f1", x"ec", x"10", x"f1", x"ef", x"13", x"08", x"25",
    x"08", x"28", x"0b", x"0d", x"f7", x"ea", x"30", x"f2",
    x"ed", x"19", x"30", x"22", x"ef", x"16", x"0b", x"fa",
    x"f4", x"ff", x"17", x"20", x"3e", x"28", x"1a", x"0a",
    x"df", x"d1", x"e9", x"fb", x"fb", x"fe", x"05", x"05",
    x"01", x"01", x"00", x"00", x"07", x"c6", x"c9", x"d7",
    x"bb", x"ea", x"0e", x"0c", x"05", x"fd", x"21", x"25",
    x"63", x"4f", x"4b", x"31", x"11", x"10", x"cc", x"ec",
    x"fd", x"df", x"e2", x"d3", x"f1", x"ec", x"01", x"cc",
    x"a5", x"cd", x"ef", x"bf", x"ba", x"10", x"a0", x"74",
    x"3e", x"f9", x"d8", x"3b", x"11", x"da", x"dc", x"04",
    x"12", x"03", x"0c", x"10", x"11", x"01", x"f4", x"e5",
    x"e7", x"e3", x"de", x"e0", x"ff", x"24", x"0d", x"f4",
    x"e5", x"e9", x"ce", x"54", x"15", x"00", x"0a", x"e2",
    x"0f", x"f0", x"de", x"b4", x"f9", x"0f", x"00", x"00",
    x"04", x"0b", x"fd", x"07", x"15", x"0c", x"17", x"1b",
    x"fd", x"1d", x"1a", x"15", x"10", x"d4", x"1d", x"f4",
    x"fc", x"3c", x"f1", x"03", x"78", x"ff", x"fa", x"fb",
    x"1d", x"3b", x"d3", x"13", x"1c", x"18", x"30", x"1b",
    x"ff", x"02", x"01", x"02", x"05", x"03", x"02", x"00",
    x"02", x"dd", x"b8", x"f5", x"e9", x"f0", x"15", x"cd",
    x"af", x"99", x"19", x"d2", x"f9", x"20", x"e0", x"d7",
    x"11", x"c7", x"7a", x"ed", x"04", x"ff", x"06", x"dd",
    x"ec", x"21", x"b5", x"ac", x"07", x"1f", x"fc", x"0c",
    x"28", x"1b", x"cd", x"01", x"14", x"19", x"f8", x"cf",
    x"eb", x"e0", x"eb", x"f6", x"f0", x"f3", x"d6", x"0b",
    x"12", x"f4", x"e2", x"04", x"0f", x"0f", x"1e", x"4a",
    x"3c", x"17", x"22", x"f7", x"f2", x"ee", x"a9", x"b7",
    x"04", x"04", x"fe", x"05", x"00", x"04", x"ff", x"fd",
    x"02", x"01", x"fd", x"fd", x"fe", x"fb", x"fd", x"04",
    x"03", x"04", x"28", x"04", x"21", x"21", x"e7", x"eb",
    x"2a", x"0a", x"3a", x"4a", x"e1", x"d6", x"e2", x"04",
    x"23", x"f8", x"02", x"2a", x"e8", x"00", x"04", x"27",
    x"30", x"fb", x"ed", x"18", x"04", x"02", x"f2", x"f7",
    x"fa", x"fb", x"f9", x"7f", x"b7", x"df", x"08", x"00",
    x"40", x"27", x"0b", x"0e", x"f7", x"ed", x"0e", x"d6",
    x"19", x"0c", x"0a", x"26", x"1e", x"39", x"1c", x"db",
    x"10", x"09", x"16", x"13", x"01", x"11", x"3d", x"d1",
    x"03", x"06", x"fe", x"0b", x"d6", x"10", x"1a", x"fa",
    x"07", x"10", x"1c", x"fc", x"f3", x"11", x"07", x"26",
    x"29", x"42", x"16", x"09", x"ef", x"11", x"c3", x"dc",
    x"a7", x"dc", x"a9", x"ac", x"09", x"22", x"13", x"05",
    x"e4", x"f5", x"05", x"f8", x"af", x"e3", x"27", x"ff",
    x"19", x"1a", x"0b", x"2c", x"0e", x"d5", x"42", x"00",
    x"de", x"41", x"ee", x"b8", x"2a", x"d3", x"ce", x"e8",
    x"ca", x"04", x"ee", x"dd", x"d6", x"13", x"e0", x"fa",
    x"ff", x"27", x"42", x"14", x"17", x"00", x"1d", x"05",
    x"f2", x"1d", x"e8", x"bc", x"e4", x"03", x"fe", x"08",
    x"46", x"0b", x"2b", x"1c", x"0f", x"04", x"2d", x"20",
    x"06", x"fa", x"05", x"0d", x"0b", x"df", x"2a", x"fa",
    x"fe", x"ca", x"fe", x"e1", x"da", x"ad", x"62", x"0a",
    x"f7", x"00", x"e6", x"0d", x"0e", x"07", x"a6", x"ce",
    x"0f", x"44", x"26", x"0c", x"46", x"f8", x"94", x"fe",
    x"13", x"cf", x"dd", x"0e", x"f1", x"fd", x"41", x"c2",
    x"06", x"25", x"0c", x"34", x"fe", x"14", x"22", x"09",
    x"e8", x"df", x"c4", x"cb", x"df", x"b8", x"08", x"c9",
    x"a2", x"d7", x"d5", x"c4", x"1b", x"c9", x"f1", x"64",
    x"e7", x"0f", x"10", x"eb", x"08", x"ea", x"ef", x"01",
    x"35", x"29", x"39", x"13", x"22", x"03", x"ff", x"1a",
    x"10", x"36", x"ed", x"ba", x"16", x"ff", x"f4", x"25",
    x"31", x"0b", x"12", x"27", x"07", x"36", x"ef", x"d2",
    x"1b", x"fe", x"91", x"23", x"38", x"5c", x"1c", x"11",
    x"f1", x"ef", x"10", x"21", x"f6", x"10", x"31", x"3f",
    x"2b", x"03", x"27", x"44", x"27", x"65", x"2f", x"fd",
    x"d8", x"10", x"f0", x"17", x"0f", x"09", x"15", x"fc",
    x"e9", x"ff", x"04", x"fb", x"fc", x"ff", x"fb", x"06",
    x"fd", x"ff", x"12", x"0f", x"21", x"13", x"13", x"18",
    x"0a", x"14", x"10", x"e2", x"e3", x"b0", x"f0", x"e1",
    x"db", x"d4", x"fd", x"3d", x"f1", x"0a", x"e5", x"e9",
    x"fe", x"ac", x"d8", x"fc", x"18", x"d3", x"c7", x"e2",
    x"fa", x"af", x"c7", x"1d", x"bf", x"a7", x"e4", x"f5",
    x"f4", x"06", x"13", x"30", x"2e", x"22", x"3d", x"c8",
    x"ab", x"61", x"d4", x"cf", x"dd", x"e7", x"d0", x"01",
    x"17", x"f8", x"00", x"33", x"17", x"00", x"e6", x"f7",
    x"22", x"23", x"3b", x"d0", x"40", x"06", x"f3", x"fb",
    x"44", x"2b", x"f6", x"ca", x"c2", x"d1", x"b4", x"b4",
    x"0d", x"04", x"d7", x"01", x"03", x"03", x"08", x"fd",
    x"ff", x"fe", x"fc", x"02", x"e6", x"dc", x"f2", x"cf",
    x"da", x"f3", x"ff", x"f0", x"ee", x"04", x"a9", x"34",
    x"e3", x"c8", x"fc", x"1b", x"cc", x"d4", x"33", x"1c",
    x"d7", x"31", x"27", x"14", x"55", x"38", x"26", x"f4",
    x"f9", x"dc", x"ca", x"e5", x"ee", x"cc", x"00", x"fa",
    x"f5", x"37", x"6a", x"ea", x"f2", x"2b", x"eb", x"f4",
    x"14", x"15", x"dd", x"1a", x"f6", x"87", x"cb", x"45",
    x"f0", x"1b", x"0c", x"60", x"42", x"04", x"3d", x"3e",
    x"27", x"58", x"3a", x"fa", x"3d", x"fd", x"26", x"f8",
    x"c7", x"05", x"e5", x"ca", x"01", x"01", x"08", x"ff",
    x"ff", x"05", x"04", x"02", x"08", x"17", x"e7", x"8b",
    x"26", x"dc", x"89", x"1c", x"d7", x"bd", x"0a", x"1c",
    x"11", x"28", x"f3", x"fe", x"2d", x"f4", x"fb", x"a3",
    x"08", x"cd", x"c4", x"0b", x"0b", x"f1", x"eb", x"09",
    x"ff", x"fc", x"fe", x"fe", x"fc", x"01", x"ff", x"fd",
    x"03", x"1e", x"0a", x"d3", x"49", x"04", x"e0", x"55",
    x"0a", x"f1", x"d5", x"bf", x"d9", x"d0", x"c6", x"c9",
    x"00", x"b5", x"76", x"fa", x"fc", x"e2", x"34", x"ec",
    x"c8", x"28", x"ff", x"e4", x"78", x"8b", x"2b", x"2c",
    x"1d", x"ed", x"2a", x"29", x"fe", x"ba", x"c9", x"e1",
    x"b9", x"a8", x"ac", x"dd", x"b6", x"97", x"0c", x"c5",
    x"22", x"0b", x"b9", x"28", x"29", x"0f", x"01", x"f0",
    x"fd", x"02", x"2b", x"20", x"3d", x"11", x"31", x"27",
    x"01", x"02", x"00", x"fb", x"01", x"ff", x"fe", x"01",
    x"07", x"03", x"fe", x"fe", x"f9", x"09", x"fc", x"02",
    x"01", x"01", x"c0", x"ca", x"c1", x"e8", x"b3", x"f5",
    x"b7", x"ba", x"e5", x"9d", x"df", x"16", x"ec", x"f8",
    x"f2", x"e8", x"07", x"1e", x"fc", x"c9", x"dc", x"14",
    x"ed", x"df", x"1d", x"54", x"17", x"f3", x"f2", x"e3",
    x"fb", x"04", x"de", x"22", x"ec", x"e0", x"16", x"28",
    x"07", x"f7", x"ff", x"13", x"16", x"fc", x"1b", x"d8",
    x"0f", x"1a", x"3a", x"30", x"1c", x"05", x"10", x"1e",
    x"15", x"f9", x"33", x"16", x"f0", x"f6", x"00", x"0e",
    x"01", x"36", x"00", x"e0", x"02", x"e6", x"07", x"0d",
    x"17", x"0c", x"e6", x"02", x"11", x"1d", x"f7", x"34",
    x"ed", x"f9", x"30", x"16", x"12", x"dd", x"32", x"33",
    x"38", x"72", x"60", x"24", x"44", x"27", x"05", x"1e",
    x"0b", x"c8", x"07", x"c5", x"b8", x"a3", x"d3", x"f6",
    x"ba", x"01", x"14", x"ec", x"2a", x"08", x"18", x"fe",
    x"e4", x"1f", x"3c", x"25", x"f9", x"45", x"fe", x"f5",
    x"3a", x"3d", x"0e", x"25", x"32", x"d8", x"34", x"15",
    x"02", x"04", x"5d", x"03", x"ca", x"a1", x"8a", x"6e",
    x"66", x"27", x"f7", x"f6", x"3d", x"ee", x"e7", x"0c",
    x"cf", x"ca", x"b7", x"ce", x"d3", x"dc", x"bc", x"be",
    x"e1", x"ae", x"b5", x"d4", x"e8", x"ff", x"0d", x"41",
    x"11", x"17", x"27", x"0e", x"e9", x"0a", x"20", x"cc",
    x"12", x"0b", x"e7", x"35", x"6c", x"ed", x"e9", x"01",
    x"f7", x"a8", x"a6", x"e9", x"cd", x"80", x"0c", x"f4",
    x"10", x"e3", x"00", x"3d", x"12", x"15", x"03", x"23",
    x"39", x"ff", x"2f", x"40", x"f6", x"b3", x"bc", x"d6",
    x"10", x"18", x"2f", x"09", x"15", x"fd", x"db", x"dc",
    x"d0", x"e7", x"e8", x"d7", x"44", x"1d", x"c4", x"2b",
    x"1a", x"3b", x"13", x"01", x"ea", x"9b", x"1a", x"1f",
    x"ff", x"86", x"1f", x"32", x"0e", x"fa", x"00", x"03",
    x"f7", x"97", x"fe", x"0a", x"ed", x"d6", x"ea", x"fb",
    x"e7", x"fa", x"1f", x"e9", x"da", x"25", x"0e", x"b9",
    x"24", x"20", x"f3", x"ed", x"07", x"54", x"00", x"1d",
    x"a8", x"3e", x"21", x"20", x"00", x"fb", x"05", x"df",
    x"03", x"f8", x"2e", x"17", x"f3", x"0c", x"c7", x"d6",
    x"04", x"24", x"24", x"ed", x"19", x"e4", x"d6", x"aa",
    x"d0", x"05", x"04", x"01", x"05", x"fd", x"03", x"ff",
    x"fd", x"04", x"fb", x"0b", x"ee", x"00", x"17", x"25",
    x"b1", x"d2", x"c2", x"14", x"fc", x"e8", x"03", x"e5",
    x"d2", x"0b", x"0c", x"1b", x"fb", x"21", x"06", x"25",
    x"25", x"2a", x"eb", x"e9", x"1d", x"d4", x"e4", x"e5",
    x"ea", x"f1", x"22", x"a7", x"f5", x"df", x"1c", x"0a",
    x"e5", x"fe", x"f0", x"be", x"cd", x"c1", x"4d", x"13",
    x"fa", x"f9", x"29", x"e9", x"e8", x"15", x"03", x"17",
    x"f2", x"4a", x"02", x"dd", x"fe", x"10", x"b6", x"b7",
    x"e8", x"2a", x"04", x"fc", x"d1", x"11", x"18", x"cc",
    x"bc", x"0c", x"1e", x"11", x"fc", x"d5", x"fe", x"f2",
    x"ab", x"b9", x"ec", x"00", x"fe", x"01", x"0b", x"03",
    x"ff", x"0c", x"06", x"00", x"4a", x"28", x"09", x"19",
    x"39", x"21", x"1c", x"17", x"0b", x"08", x"16", x"ea",
    x"b5", x"eb", x"ea", x"2a", x"22", x"55", x"13", x"05",
    x"d5", x"45", x"57", x"57", x"45", x"1c", x"58", x"0d",
    x"f4", x"2e", x"20", x"10", x"01", x"d3", x"da", x"ba",
    x"d7", x"f1", x"0c", x"fd", x"f3", x"1f", x"ef", x"17",
    x"3f", x"df", x"f4", x"11", x"4e", x"2f", x"ea", x"16",
    x"e4", x"f2", x"ee", x"04", x"10", x"09", x"0c", x"19",
    x"f1", x"b7", x"71", x"ff", x"07", x"26", x"07", x"f0",
    x"e5", x"92", x"19", x"1f", x"09", x"0e", x"0d", x"12",
    x"0e", x"08", x"0b", x"10", x"0b", x"07", x"10", x"fe",
    x"03", x"0f", x"25", x"2c", x"4d", x"4a", x"d1", x"ee",
    x"f3", x"0f", x"f0", x"e4", x"d5", x"eb", x"d6", x"0c",
    x"f9", x"fd", x"e7", x"e9", x"fd", x"da", x"fa", x"02",
    x"ff", x"fd", x"01", x"03", x"05", x"fe", x"01", x"fd",
    x"fc", x"54", x"29", x"23", x"3d", x"1f", x"f5", x"dc",
    x"09", x"26", x"3c", x"36", x"37", x"48", x"08", x"fd",
    x"fd", x"15", x"f4", x"12", x"f9", x"dc", x"f6", x"0d",
    x"01", x"b8", x"e9", x"ef", x"fb", x"09", x"ea", x"e0",
    x"f1", x"e3", x"db", x"21", x"33", x"da", x"d2", x"04",
    x"17", x"11", x"d6", x"bd", x"c1", x"b0", x"08", x"d5",
    x"ff", x"e3", x"f1", x"d5", x"1b", x"1c", x"02", x"d9",
    x"c3", x"ec", x"0b", x"09", x"d4", x"dd", x"09", x"dd",
    x"fa", x"04", x"ff", x"07", x"07", x"01", x"01", x"04",
    x"00", x"f9", x"01", x"fe", x"ff", x"08", x"fb", x"02",
    x"01", x"fe", x"cd", x"f5", x"dd", x"97", x"98", x"8d",
    x"9b", x"b6", x"93", x"d5", x"f2", x"d6", x"fb", x"12",
    x"27", x"dd", x"0a", x"12", x"fb", x"f0", x"cb", x"dd",
    x"0d", x"ea", x"09", x"36", x"1b", x"24", x"20", x"12",
    x"f9", x"d5", x"cf", x"3f", x"bf", x"da", x"11", x"eb",
    x"0a", x"bb", x"b7", x"a0", x"f6", x"dd", x"f9", x"eb",
    x"e9", x"ea", x"c3", x"27", x"34", x"d1", x"eb", x"f8",
    x"fa", x"25", x"f9", x"e7", x"fe", x"28", x"5b", x"3c",
    x"35", x"33", x"d6", x"10", x"dd", x"d6", x"e2", x"fc",
    x"ed", x"bf", x"c6", x"06", x"2f", x"e6", x"ec", x"08",
    x"dc", x"d2", x"dd", x"0f", x"05", x"0b", x"02", x"f5",
    x"24", x"8d", x"a6", x"cd", x"5b", x"40", x"30", x"14",
    x"b5", x"7c", x"fe", x"f2", x"f7", x"0c", x"31", x"0e",
    x"1c", x"19", x"f3", x"f7", x"0d", x"44", x"2c", x"37",
    x"35", x"19", x"44", x"2c", x"24", x"e8", x"f6", x"eb",
    x"06", x"30", x"e1", x"cd", x"04", x"e6", x"20", x"e0",
    x"18", x"f9", x"2f", x"ff", x"f5", x"f9", x"14", x"da",
    x"0c", x"67", x"2e", x"3d", x"79", x"20", x"02", x"35",
    x"1b", x"01", x"01", x"2c", x"f9", x"fb", x"02", x"f4",
    x"0e", x"16", x"0c", x"d2", x"b7", x"bb", x"a8", x"db",
    x"df", x"d1", x"af", x"d1", x"3e", x"2d", x"56", x"36",
    x"2d", x"53", x"23", x"30", x"22", x"ed", x"0c", x"2a",
    x"0b", x"de", x"f1", x"e8", x"e0", x"bc", x"e1", x"c0",
    x"bc", x"fb", x"bb", x"99", x"b0", x"aa", x"dc", x"4c",
    x"33", x"53", x"22", x"2c", x"18", x"2c", x"25", x"3c",
    x"26", x"11", x"2d", x"11", x"10", x"10", x"14", x"08",
    x"0c", x"fb", x"0d", x"04", x"1c", x"1b", x"1f", x"1c",
    x"33", x"39", x"d1", x"11", x"06", x"ab", x"08", x"06",
    x"ff", x"4d", x"16", x"e8", x"da", x"09", x"be", x"d6",
    x"f6", x"1d", x"07", x"12", x"18", x"19", x"0e", x"17",
    x"25", x"1a", x"f9", x"18", x"f5", x"f5", x"03", x"39",
    x"f8", x"f1", x"23", x"10", x"e6", x"2d", x"15", x"f2",
    x"0b", x"de", x"f0", x"fd", x"08", x"e2", x"cc", x"f8",
    x"d0", x"c8", x"f4", x"f8", x"17", x"01", x"01", x"07",
    x"0d", x"26", x"60", x"eb", x"1f", x"3b", x"e0", x"d9",
    x"0d", x"03", x"fe", x"fc", x"fb", x"02", x"fd", x"01",
    x"fe", x"04", x"03", x"0d", x"07", x"c6", x"d4", x"03",
    x"e1", x"ec", x"02", x"e3", x"fe", x"05", x"19", x"0a",
    x"f7", x"2a", x"4a", x"ce", x"e2", x"15", x"1f", x"25",
    x"4e", x"2e", x"49", x"47", x"21", x"03", x"e5", x"fd",
    x"fd", x"00", x"12", x"15", x"33", x"27", x"19", x"03",
    x"c5", x"12", x"cc", x"d4", x"19", x"d0", x"9e", x"06",
    x"18", x"1c", x"1e", x"18", x"06", x"1d", x"02", x"35",
    x"0a", x"2f", x"17", x"32", x"03", x"fe", x"4d", x"cd",
    x"02", x"bd", x"10", x"0e", x"d4", x"f2", x"e2", x"2d",
    x"ef", x"ec", x"02", x"33", x"2e", x"1e", x"23", x"15",
    x"6d", x"2e", x"fe", x"ff", x"00", x"fe", x"f9", x"fb",
    x"fc", x"07", x"05", x"fc", x"39", x"4a", x"30", x"19",
    x"34", x"48", x"1e", x"27", x"3e", x"13", x"fe", x"e0",
    x"1c", x"1e", x"01", x"09", x"fb", x"20", x"f2", x"eb",
    x"2c", x"f6", x"f8", x"2a", x"f7", x"0f", x"25", x"1f",
    x"31", x"1e", x"2d", x"1f", x"12", x"2a", x"2c", x"3c",
    x"44", x"df", x"ea", x"e1", x"df", x"f5", x"06", x"e4",
    x"e5", x"f9", x"33", x"2e", x"2f", x"02", x"11", x"14",
    x"f1", x"f8", x"2c", x"00", x"ec", x"07", x"e6", x"e9",
    x"eb", x"e2", x"f5", x"fb", x"19", x"ff", x"e0", x"26",
    x"17", x"2e", x"2d", x"29", x"0e", x"08", x"05", x"05",
    x"01", x"05", x"03", x"02", x"0d", x"59", x"33", x"2b",
    x"f5", x"2b", x"24", x"e1", x"3b", x"46", x"f3", x"2a",
    x"f1", x"da", x"db", x"f1", x"e5", x"dc", x"e0", x"01",
    x"ec", x"18", x"d9", x"ef", x"ce", x"1a", x"e5", x"d6",
    x"01", x"01", x"fe", x"ff", x"03", x"05", x"fb", x"ff",
    x"00", x"c9", x"e0", x"17", x"f9", x"02", x"18", x"ff",
    x"fe", x"10", x"28", x"60", x"32", x"20", x"2d", x"4c",
    x"46", x"39", x"4b", x"f7", x"f6", x"04", x"f3", x"05",
    x"14", x"ff", x"21", x"0e", x"15", x"06", x"2e", x"f8",
    x"09", x"21", x"b7", x"c6", x"e1", x"a1", x"8e", x"87",
    x"69", x"5f", x"42", x"52", x"3d", x"ec", x"22", x"09",
    x"2e", x"d3", x"c5", x"ea", x"f0", x"fa", x"02", x"df",
    x"b5", x"0b", x"f2", x"bf", x"cc", x"e4", x"dd", x"ae",
    x"02", x"fc", x"00", x"f4", x"fb", x"01", x"03", x"fe",
    x"00", x"f9", x"f8", x"fc", x"00", x"fb", x"fa", x"01",
    x"fb", x"ff", x"fd", x"0a", x"08", x"ff", x"f7", x"0a",
    x"f9", x"02", x"01", x"f2", x"dd", x"11", x"f1", x"ec",
    x"e9", x"08", x"ee", x"e3", x"f7", x"00", x"fa", x"1a",
    x"0a", x"e6", x"07", x"f1", x"e6", x"20", x"f5", x"fa",
    x"f7", x"d3", x"fa", x"e4", x"fd", x"13", x"dc", x"af",
    x"e2", x"e3", x"c6", x"04", x"ed", x"e5", x"df", x"49",
    x"f0", x"df", x"38", x"11", x"ca", x"ee", x"aa", x"cf",
    x"0f", x"e1", x"e4", x"2a", x"b8", x"ff", x"80", x"19",
    x"2e", x"4c", x"14", x"1e", x"38", x"37", x"16", x"3b",
    x"43", x"22", x"bf", x"d0", x"cc", x"fa", x"f6", x"f1",
    x"13", x"da", x"d3", x"fd", x"de", x"06", x"f1", x"0f",
    x"0b", x"08", x"07", x"f2", x"25", x"2f", x"52", x"43",
    x"51", x"4a", x"4e", x"5b", x"62", x"34", x"2f", x"15",
    x"0c", x"07", x"10", x"17", x"23", x"1a", x"1c", x"f4",
    x"d8", x"05", x"d9", x"08", x"fe", x"0a", x"fd", x"0b",
    x"e9", x"e3", x"f3", x"eb", x"e4", x"12", x"b3", x"ad",
    x"db", x"fb", x"78", x"b5", x"df", x"03", x"c4", x"d2",
    x"91", x"dc", x"c8", x"b1", x"16", x"05", x"01", x"04",
    x"0f", x"d3", x"22", x"35", x"21", x"15", x"0f", x"1b",
    x"24", x"20", x"1d", x"23", x"1b", x"d9", x"02", x"f6",
    x"c5", x"f4", x"0f", x"ff", x"0e", x"2f", x"fc", x"c1",
    x"e8", x"f0", x"6f", x"e4", x"05", x"e3", x"e4", x"ea",
    x"e6", x"04", x"ff", x"fc", x"02", x"f7", x"10", x"17",
    x"23", x"d8", x"16", x"38", x"34", x"4c", x"4a", x"f5",
    x"fb", x"c6", x"e0", x"ce", x"a4", x"bc", x"ab", x"c9",
    x"c1", x"d7", x"fd", x"e1", x"c5", x"0d", x"bf", x"d5",
    x"11", x"d9", x"dd", x"08", x"18", x"26", x"19", x"54",
    x"11", x"03", x"02", x"1f", x"29", x"2c", x"c1", x"f4",
    x"05", x"cc", x"a9", x"1b", x"0d", x"ff", x"6f", x"07",
    x"f7", x"35", x"db", x"00", x"21", x"af", x"cd", x"db",
    x"03", x"20", x"25", x"0b", x"09", x"34", x"21", x"01",
    x"0e", x"2c", x"17", x"fa", x"da", x"c8", x"05", x"f6",
    x"ec", x"04", x"22", x"01", x"e6", x"38", x"36", x"2d",
    x"2d", x"01", x"14", x"0e", x"06", x"36", x"22", x"ca",
    x"cb", x"88", x"8e", x"07", x"ce", x"e1", x"1f", x"fb",
    x"01", x"fb", x"01", x"fc", x"04", x"fe", x"04", x"06",
    x"fb", x"00", x"90", x"da", x"03", x"f7", x"eb", x"f2",
    x"e3", x"d9", x"f3", x"18", x"27", x"07", x"2e", x"26",
    x"cf", x"0f", x"e6", x"db", x"eb", x"0a", x"37", x"34",
    x"34", x"24", x"0b", x"2f", x"f6", x"01", x"1e", x"29",
    x"b8", x"10", x"30", x"e0", x"e3", x"e7", x"a3", x"ce",
    x"e8", x"ab", x"df", x"1f", x"e4", x"e1", x"e8", x"1d",
    x"c1", x"df", x"dc", x"b2", x"ea", x"dd", x"ee", x"c8",
    x"dc", x"e5", x"2e", x"28", x"fd", x"17", x"55", x"f4",
    x"ff", x"25", x"1a", x"07", x"04", x"e3", x"de", x"e2",
    x"d7", x"e5", x"0e", x"f9", x"22", x"a6", x"c1", x"f0",
    x"0a", x"de", x"b8", x"ff", x"02", x"ff", x"00", x"fe",
    x"fb", x"00", x"03", x"fc", x"df", x"dd", x"ea", x"cf",
    x"e9", x"03", x"d6", x"e1", x"f3", x"ba", x"86", x"0a",
    x"ac", x"f9", x"15", x"7b", x"3d", x"1e", x"3c", x"43",
    x"fc", x"1a", x"25", x"16", x"f5", x"16", x"06", x"04",
    x"d2", x"d8", x"04", x"da", x"d9", x"fa", x"fa", x"dc",
    x"cf", x"bc", x"30", x"e5", x"dd", x"19", x"f4", x"cd",
    x"db", x"d3", x"f6", x"0e", x"ee", x"fa", x"f4", x"19",
    x"1b", x"b2", x"e5", x"f9", x"e0", x"01", x"e6", x"d1",
    x"e7", x"ba", x"c5", x"cd", x"e5", x"ed", x"ba", x"32",
    x"fa", x"d6", x"fe", x"f2", x"05", x"0c", x"0b", x"08",
    x"0d", x"07", x"03", x"08", x"fd", x"d8", x"d3", x"e8",
    x"ab", x"c6", x"d8", x"f8", x"01", x"00", x"e6", x"0a",
    x"12", x"fc", x"30", x"2e", x"f4", x"02", x"13", x"f2",
    x"35", x"3c", x"fc", x"17", x"00", x"ed", x"f5", x"0b",
    x"fc", x"05", x"ff", x"fa", x"00", x"02", x"fd", x"ff",
    x"02", x"21", x"67", x"58", x"1e", x"1e", x"01", x"0a",
    x"15", x"0e", x"f6", x"2c", x"4d", x"f6", x"16", x"1e",
    x"e2", x"c7", x"ab", x"25", x"48", x"3a", x"d2", x"05",
    x"f9", x"37", x"1e", x"07", x"c4", x"b5", x"bc", x"e2",
    x"a9", x"e5", x"1b", x"0d", x"10", x"bd", x"d1", x"e4",
    x"0c", x"f4", x"14", x"f7", x"fc", x"00", x"e2", x"c7",
    x"e6", x"04", x"f0", x"13", x"07", x"14", x"0a", x"40",
    x"25", x"3d", x"02", x"fd", x"47", x"06", x"df", x"06",
    x"fd", x"00", x"05", x"03", x"01", x"fe", x"fe", x"00",
    x"05", x"fd", x"fc", x"01", x"fe", x"01", x"00", x"fe",
    x"fe", x"03", x"c6", x"d2", x"af", x"d2", x"e9", x"ea",
    x"a0", x"d4", x"df", x"c7", x"cc", x"13", x"e9", x"f7",
    x"00", x"dd", x"dd", x"ec", x"1b", x"fa", x"fe", x"d7",
    x"e3", x"dc", x"00", x"13", x"d9", x"e9", x"09", x"d2",
    x"38", x"2f", x"f7", x"f1", x"87", x"c9", x"eb", x"ce",
    x"06", x"b5", x"e1", x"f6", x"d3", x"c5", x"e0", x"2a",
    x"e4", x"0e", x"f7", x"1b", x"17", x"2d", x"4d", x"13",
    x"ca", x"f4", x"4b", x"73", x"e8", x"1d", x"e5", x"cf",
    x"ff", x"0b", x"21", x"db", x"3f", x"0d", x"f7", x"00",
    x"fc", x"08", x"d0", x"23", x"0c", x"e7", x"0a", x"11",
    x"5c", x"28", x"32", x"01", x"f3", x"ea", x"f2", x"c8",
    x"b1", x"9b", x"ce", x"0e", x"e4", x"f6", x"05", x"19",
    x"07", x"fd", x"11", x"11", x"ff", x"10", x"15", x"f3",
    x"f3", x"0b", x"15", x"30", x"30", x"2d", x"c9", x"f9",
    x"eb", x"dd", x"eb", x"0c", x"0d", x"d2", x"b1", x"d9",
    x"87", x"8b", x"f7", x"d3", x"b3", x"1e", x"ff", x"14",
    x"df", x"36", x"fc", x"c6", x"1c", x"2b", x"c8", x"e5",
    x"41", x"eb", x"0d", x"24", x"09", x"0a", x"09", x"03",
    x"1c", x"1a", x"ac", x"ea", x"eb", x"cc", x"d2", x"19",
    x"de", x"ce", x"e9", x"1e", x"10", x"02", x"08", x"f6",
    x"11", x"04", x"fe", x"07", x"11", x"ff", x"1b", x"de",
    x"04", x"fa", x"fa", x"e3", x"e9", x"a1", x"09", x"30",
    x"cc", x"f2", x"1b", x"d0", x"8a", x"a8", x"28", x"fa",
    x"15", x"11", x"08", x"13", x"2e", x"10", x"20", x"52",
    x"8e", x"34", x"26", x"2f", x"d8", x"15", x"1f", x"c0",
    x"ff", x"36", x"63", x"0c", x"10", x"17", x"d4", x"e0",
    x"19", x"0b", x"e0", x"0d", x"34", x"19", x"08", x"50",
    x"56", x"1e", x"b2", x"09", x"1d", x"a3", x"df", x"f2",
    x"27", x"8e", x"2e", x"fe", x"eb", x"dd", x"28", x"1d",
    x"0b", x"33", x"1b", x"f9", x"0c", x"de", x"eb", x"ae",
    x"a3", x"b2", x"e2", x"ab", x"d1", x"c8", x"cf", x"8c",
    x"0b", x"fa", x"d8", x"1d", x"32", x"fc", x"0b", x"f8",
    x"dc", x"33", x"26", x"08", x"10", x"3b", x"10", x"19",
    x"ec", x"11", x"37", x"6b", x"34", x"26", x"2b", x"e4",
    x"18", x"19", x"38", x"16", x"43", x"27", x"f3", x"cf",
    x"d5", x"01", x"03", x"fb", x"01", x"fc", x"fc", x"fd",
    x"fb", x"fc", x"e4", x"1a", x"df", x"56", x"31", x"23",
    x"cc", x"f7", x"e8", x"be", x"e7", x"06", x"ed", x"eb",
    x"fa", x"0a", x"09", x"cf", x"c0", x"ac", x"77", x"12",
    x"0a", x"ba", x"32", x"42", x"14", x"bd", x"e2", x"de",
    x"cb", x"de", x"eb", x"cd", x"e3", x"db", x"f1", x"ed",
    x"0e", x"12", x"04", x"15", x"0d", x"ea", x"da", x"ed",
    x"f5", x"0e", x"fe", x"04", x"07", x"fe", x"da", x"e5",
    x"06", x"fc", x"f8", x"b9", x"4d", x"35", x"fa", x"e8",
    x"00", x"e3", x"e1", x"ee", x"e4", x"ee", x"f7", x"ba",
    x"11", x"2f", x"b2", x"ea", x"e8", x"15", x"01", x"e4",
    x"6e", x"ce", x"cd", x"fa", x"01", x"fc", x"05", x"00",
    x"f7", x"ff", x"03", x"f8", x"46", x"64", x"38", x"2e",
    x"15", x"05", x"2c", x"3a", x"2b", x"e2", x"f2", x"21",
    x"e5", x"02", x"50", x"d2", x"f2", x"e5", x"03", x"f6",
    x"ca", x"42", x"28", x"17", x"3c", x"53", x"62", x"10",
    x"06", x"32", x"3a", x"2b", x"34", x"fd", x"10", x"1e",
    x"e0", x"04", x"f2", x"cc", x"e9", x"c9", x"d3", x"ea",
    x"d7", x"d5", x"d7", x"f4", x"24", x"0d", x"fd", x"21",
    x"2e", x"c8", x"e2", x"e9", x"d1", x"c3", x"14", x"18",
    x"fc", x"f8", x"05", x"e8", x"0d", x"31", x"0d", x"ff",
    x"fa", x"d5", x"05", x"02", x"00", x"ff", x"03", x"0b",
    x"fc", x"00", x"07", x"07", x"02", x"d4", x"e5", x"c7",
    x"06", x"f5", x"f6", x"29", x"f3", x"fd", x"1c", x"47",
    x"22", x"eb", x"31", x"16", x"d8", x"13", x"08", x"2e",
    x"08", x"21", x"14", x"33", x"32", x"ec", x"0e", x"14",
    x"01", x"00", x"04", x"00", x"ff", x"fd", x"fc", x"ff",
    x"06", x"1e", x"15", x"f5", x"20", x"14", x"23", x"10",
    x"0b", x"16", x"61", x"2a", x"11", x"2f", x"0d", x"10",
    x"09", x"e9", x"1b", x"d1", x"12", x"f7", x"fc", x"0b",
    x"0c", x"0b", x"24", x"0a", x"28", x"e6", x"26", x"ec",
    x"ab", x"a0", x"c7", x"ac", x"b0", x"f2", x"c5", x"0b",
    x"f7", x"dd", x"df", x"d3", x"e9", x"19", x"d7", x"cc",
    x"0e", x"ec", x"c2", x"0e", x"05", x"18", x"e6", x"d7",
    x"df", x"ec", x"e0", x"f2", x"ed", x"f1", x"ea", x"b0",
    x"00", x"01", x"02", x"fd", x"01", x"fb", x"02", x"fe",
    x"07", x"fe", x"ff", x"00", x"ff", x"fe", x"fc", x"f8",
    x"03", x"02", x"fb", x"ee", x"1a", x"b2", x"c8", x"ec",
    x"90", x"95", x"a9", x"e8", x"f9", x"c8", x"e0", x"eb",
    x"cc", x"f2", x"07", x"11", x"74", x"a8", x"b3", x"e3",
    x"dc", x"cf", x"f3", x"fe", x"19", x"38", x"1b", x"1e",
    x"35", x"2a", x"df", x"b9", x"d6", x"9e", x"0d", x"13",
    x"0c", x"4c", x"f6", x"e8", x"d5", x"cb", x"a7", x"e1",
    x"e6", x"f0", x"d8", x"37", x"19", x"09", x"0e", x"28",
    x"e2", x"06", x"f7", x"e2", x"ef", x"1d", x"be", x"eb",
    x"1f", x"31", x"f1", x"df", x"e5", x"01", x"d3", x"d7",
    x"e4", x"02", x"f3", x"f5", x"fb", x"16", x"fb", x"f1",
    x"20", x"e6", x"f3", x"0b", x"e0", x"fd", x"1e", x"f6",
    x"ed", x"d0", x"05", x"0d", x"13", x"8c", x"47", x"2c",
    x"f0", x"13", x"03", x"e5", x"e7", x"d9", x"20", x"2c",
    x"05", x"0a", x"ed", x"08", x"07", x"fd", x"29", x"31",
    x"ff", x"e8", x"20", x"28", x"e7", x"f0", x"14", x"6b",
    x"d9", x"12", x"a8", x"f0", x"11", x"ab", x"cb", x"d3",
    x"22", x"cd", x"93", x"f6", x"e2", x"00", x"1a", x"1f",
    x"14", x"32", x"20", x"0e", x"ec", x"f4", x"af", x"39",
    x"29", x"12", x"f6", x"f2", x"20", x"a4", x"d0", x"fa",
    x"ac", x"f8", x"e8", x"98", x"4f", x"df", x"f9", x"b2",
    x"c7", x"05", x"1d", x"c4", x"d0", x"e6", x"00", x"24",
    x"0a", x"af", x"f1", x"25", x"16", x"1e", x"f7", x"1e",
    x"2e", x"24", x"18", x"2b", x"f5", x"dc", x"fe", x"11",
    x"ec", x"01", x"18", x"54", x"f1", x"01", x"18", x"9e",
    x"f3", x"f8", x"25", x"22", x"15", x"e5", x"fd", x"46",
    x"2a", x"fc", x"d0", x"f4", x"11", x"11", x"fa", x"e7",
    x"e6", x"0c", x"1f", x"13", x"c0", x"ca", x"ec", x"ae",
    x"c5", x"e3", x"1a", x"3b", x"30", x"0a", x"b6", x"bd",
    x"04", x"bc", x"d7", x"05", x"b7", x"ff", x"05", x"09",
    x"fa", x"3a", x"18", x"20", x"07", x"e1", x"c8", x"30",
    x"05", x"fc", x"11", x"15", x"1b", x"0d", x"10", x"4f",
    x"ed", x"e2", x"53", x"e3", x"e5", x"11", x"f4", x"e6",
    x"ff", x"c4", x"ff", x"36", x"e5", x"ea", x"f4", x"c6",
    x"e9", x"e5", x"90", x"ea", x"f6", x"ee", x"f8", x"42",
    x"2c", x"01", x"05", x"d7", x"0f", x"1c", x"20", x"d8",
    x"33", x"fb", x"fd", x"02", x"fb", x"05", x"fb", x"fb",
    x"fb", x"01", x"21", x"36", x"43", x"2c", x"f5", x"0b",
    x"f5", x"f5", x"1c", x"20", x"40", x"36", x"7d", x"db",
    x"d9", x"e2", x"eb", x"32", x"c7", x"f4", x"3c", x"3a",
    x"f4", x"0b", x"1f", x"32", x"38", x"2d", x"26", x"1c",
    x"03", x"02", x"f6", x"db", x"be", x"f9", x"28", x"0f",
    x"da", x"e4", x"fc", x"ce", x"0d", x"ff", x"0e", x"d0",
    x"27", x"12", x"49", x"f6", x"e8", x"fb", x"f6", x"d0",
    x"25", x"e7", x"ed", x"42", x"a7", x"b9", x"f0", x"c3",
    x"d1", x"26", x"28", x"38", x"12", x"d7", x"b8", x"00",
    x"41", x"de", x"61", x"2a", x"35", x"c1", x"b2", x"b8",
    x"e3", x"36", x"08", x"04", x"f5", x"00", x"f8", x"f7",
    x"f8", x"08", x"fb", x"f7", x"0d", x"36", x"1c", x"ce",
    x"fb", x"0b", x"26", x"21", x"eb", x"e2", x"49", x"1f",
    x"57", x"46", x"28", x"bf", x"2b", x"11", x"ba", x"ff",
    x"05", x"04", x"d6", x"c4", x"02", x"f9", x"01", x"f4",
    x"00", x"25", x"07", x"09", x"04", x"1b", x"17", x"0b",
    x"e9", x"b3", x"d0", x"2e", x"2d", x"f1", x"06", x"1b",
    x"1c", x"16", x"09", x"08", x"e6", x"b2", x"26", x"e8",
    x"f3", x"f3", x"e3", x"c7", x"ba", x"21", x"12", x"ba",
    x"28", x"49", x"13", x"46", x"fc", x"ff", x"0d", x"17",
    x"12", x"ff", x"19", x"db", x"09", x"0e", x"0d", x"06",
    x"0b", x"0c", x"01", x"13", x"11", x"a3", x"45", x"36",
    x"fa", x"07", x"07", x"1b", x"79", x"d2", x"57", x"ce",
    x"f6", x"e8", x"dd", x"f8", x"f6", x"f5", x"ea", x"4c",
    x"26", x"05", x"ed", x"0a", x"1f", x"98", x"f3", x"2f",
    x"03", x"02", x"ff", x"02", x"00", x"fd", x"05", x"00",
    x"ff", x"f1", x"e9", x"02", x"e4", x"dc", x"f6", x"d1",
    x"d2", x"e7", x"dc", x"db", x"11", x"27", x"fe", x"fd",
    x"d9", x"c5", x"bb", x"51", x"26", x"09", x"1e", x"b7",
    x"9a", x"58", x"7f", x"62", x"c1", x"f5", x"f6", x"f7",
    x"fe", x"32", x"f6", x"e0", x"9c", x"f2", x"02", x"2a",
    x"fa", x"0a", x"01", x"c8", x"b8", x"e0", x"09", x"21",
    x"df", x"16", x"ff", x"01", x"d5", x"05", x"2f", x"3d",
    x"07", x"23", x"23", x"00", x"16", x"ad", x"ef", x"e2",
    x"fc", x"fc", x"00", x"01", x"08", x"01", x"01", x"fd",
    x"02", x"05", x"fe", x"00", x"03", x"ff", x"02", x"fc",
    x"03", x"ff", x"13", x"37", x"30", x"00", x"e7", x"fa",
    x"7c", x"ba", x"ee", x"29", x"20", x"2b", x"35", x"1b",
    x"14", x"1c", x"0d", x"36", x"2a", x"21", x"1b", x"f3",
    x"dc", x"37", x"d6", x"db", x"29", x"da", x"f3", x"cf",
    x"01", x"ff", x"fc", x"00", x"f5", x"34", x"15", x"56",
    x"de", x"3a", x"04", x"fc", x"fa", x"e0", x"08", x"09",
    x"eb", x"e8", x"37", x"45", x"51", x"bf", x"36", x"47",
    x"22", x"0a", x"f8", x"d0", x"c5", x"f0", x"84", x"ca",
    x"f5", x"20", x"1d", x"21", x"07", x"2d", x"fa", x"1e",
    x"18", x"01", x"fd", x"e4", x"8c", x"f6", x"1d", x"3e",
    x"f1", x"1f", x"39", x"ee", x"e5", x"ff", x"04", x"e0",
    x"a8", x"e5", x"d9", x"a4", x"16", x"03", x"e3", x"fd",
    x"00", x"0b", x"f3", x"15", x"ee", x"3f", x"2e", x"20",
    x"f4", x"20", x"0a", x"c2", x"f8", x"01", x"03", x"c6",
    x"71", x"29", x"e5", x"f3", x"05", x"04", x"f8", x"0c",
    x"ed", x"ab", x"2c", x"2e", x"cd", x"f6", x"e5", x"f7",
    x"e0", x"c7", x"db", x"d8", x"d7", x"33", x"ed", x"de",
    x"91", x"fb", x"ec", x"d0", x"f4", x"e0", x"04", x"39",
    x"11", x"11", x"0b", x"11", x"29", x"17", x"27", x"35",
    x"ea", x"00", x"ba", x"a5", x"9e", x"e3", x"0b", x"11",
    x"e8", x"23", x"e9", x"e6", x"db", x"0c", x"19", x"34",
    x"52", x"5d", x"38", x"4e", x"10", x"eb", x"e4", x"00",
    x"fc", x"23", x"33", x"cd", x"39", x"02", x"2e", x"0f",
    x"fd", x"d9", x"19", x"00", x"f7", x"13", x"9f", x"48",
    x"47", x"4a", x"1c", x"ea", x"ca", x"fe", x"0a", x"03",
    x"2e", x"4f", x"5d", x"2f", x"08", x"fc", x"00", x"fe",
    x"0e", x"20", x"ff", x"e5", x"d5", x"df", x"08", x"81",
    x"b0", x"d2", x"0c", x"d4", x"b0", x"12", x"e7", x"01",
    x"fa", x"08", x"04", x"fc", x"f3", x"f0", x"d0", x"d3",
    x"ad", x"e3", x"c9", x"11", x"37", x"14", x"2f", x"d1",
    x"16", x"23", x"fd", x"14", x"f1", x"0e", x"24", x"43",
    x"1b", x"ff", x"e3", x"f4", x"e6", x"07", x"12", x"ee",
    x"36", x"ff", x"1a", x"3e", x"59", x"1b", x"c3", x"0a",
    x"47", x"20", x"38", x"f6", x"b8", x"d2", x"9e", x"fc",
    x"03", x"00", x"0d", x"0d", x"e1", x"e0", x"fd", x"0b",
    x"e2", x"03", x"03", x"01", x"fd", x"02", x"01", x"05",
    x"fc", x"fc", x"16", x"51", x"23", x"3b", x"fe", x"fa",
    x"ed", x"e0", x"03", x"0a", x"0b", x"f3", x"ee", x"da",
    x"bd", x"c9", x"d4", x"1c", x"18", x"15", x"14", x"23",
    x"de", x"a2", x"08", x"fb", x"18", x"2d", x"08", x"05",
    x"f9", x"fa", x"9f", x"7b", x"93", x"bf", x"18", x"d6",
    x"c6", x"20", x"e1", x"13", x"26", x"04", x"f1", x"ff",
    x"4c", x"3e", x"20", x"41", x"08", x"13", x"3c", x"2d",
    x"18", x"15", x"2c", x"1f", x"38", x"30", x"e0", x"47",
    x"16", x"2f", x"f6", x"e8", x"ec", x"e6", x"d8", x"e8",
    x"0d", x"30", x"44", x"1c", x"04", x"0f", x"01", x"ec",
    x"9b", x"f6", x"f7", x"fe", x"fd", x"04", x"06", x"0a",
    x"07", x"03", x"04", x"04", x"39", x"33", x"3e", x"f7",
    x"0d", x"0e", x"0d", x"f4", x"18", x"f9", x"d8", x"02",
    x"1b", x"9f", x"df", x"b3", x"96", x"f4", x"05", x"df",
    x"00", x"fc", x"f4", x"ef", x"e2", x"b2", x"dd", x"33",
    x"23", x"4f", x"2a", x"1f", x"f7", x"0a", x"f1", x"0e",
    x"00", x"28", x"03", x"08", x"0e", x"2e", x"14", x"1f",
    x"1d", x"34", x"0d", x"09", x"ff", x"e7", x"e7", x"bf",
    x"d7", x"0f", x"f3", x"de", x"0f", x"f8", x"df", x"eb",
    x"bb", x"c3", x"e6", x"27", x"45", x"1a", x"bf", x"b2",
    x"b0", x"06", x"a2", x"d4", x"fe", x"03", x"0f", x"02",
    x"03", x"08", x"03", x"07", x"10", x"e2", x"08", x"0b",
    x"f4", x"ec", x"a7", x"f7", x"ad", x"e2", x"19", x"22",
    x"12", x"0c", x"46", x"54", x"15", x"03", x"0d", x"14",
    x"2c", x"3a", x"29", x"11", x"23", x"73", x"4c", x"19",
    x"fe", x"ff", x"05", x"04", x"04", x"05", x"ff", x"02",
    x"03", x"d7", x"0e", x"30", x"c5", x"e4", x"ee", x"b6",
    x"a9", x"dd", x"25", x"e5", x"1d", x"1f", x"02", x"e5",
    x"f9", x"c9", x"e3", x"31", x"d0", x"cd", x"02", x"d3",
    x"01", x"0f", x"16", x"2d", x"38", x"33", x"20", x"1f",
    x"2a", x"17", x"25", x"01", x"01", x"eb", x"1e", x"32",
    x"ef", x"e3", x"fb", x"2f", x"2a", x"f3", x"e3", x"b0",
    x"f1", x"ee", x"c6", x"e4", x"e7", x"bd", x"dd", x"2c",
    x"46", x"e7", x"0a", x"05", x"37", x"e4", x"3b", x"23",
    x"01", x"00", x"fc", x"fd", x"f7", x"fb", x"05", x"fa",
    x"fe", x"fa", x"fc", x"f7", x"03", x"fe", x"01", x"01",
    x"f9", x"03", x"db", x"f4", x"e1", x"26", x"22", x"47",
    x"12", x"1a", x"10", x"15", x"08", x"2f", x"e9", x"e9",
    x"37", x"22", x"1d", x"ca", x"f4", x"ff", x"d6", x"e7",
    x"f8", x"ee", x"8e", x"92", x"c3", x"23", x"30", x"1f",
    x"03", x"de", x"d2", x"a6", x"00", x"07", x"04", x"1d",
    x"00", x"13", x"e9", x"09", x"05", x"e8", x"d2", x"12",
    x"16", x"0e", x"4d", x"27", x"2e", x"1c", x"fc", x"c6",
    x"cb", x"a9", x"18", x"98", x"c6", x"f1", x"39", x"d5",
    x"03", x"f6", x"14", x"05", x"a9", x"f7", x"09", x"ce",
    x"01", x"43", x"00", x"e9", x"25", x"02", x"19", x"35",
    x"06", x"f5", x"01", x"fe", x"0d", x"0a", x"0a", x"fe",
    x"df", x"d1", x"cf", x"c9", x"37", x"ca", x"04", x"bf",
    x"a2", x"fa", x"bf", x"c8", x"e0", x"1a", x"05", x"e4",
    x"07", x"cd", x"de", x"96", x"f1", x"1d", x"09", x"11",
    x"12", x"10", x"f7", x"30", x"ee", x"03", x"29", x"e2",
    x"f5", x"39", x"28", x"06", x"2f", x"09", x"06", x"f1",
    x"01", x"fc", x"02", x"fb", x"fd", x"01", x"fe", x"fb",
    x"fc", x"01", x"fd", x"fb", x"00", x"fe", x"f8", x"fc",
    x"fa", x"fe", x"01", x"ff", x"fc", x"01", x"fa", x"01",
    x"02", x"00", x"07", x"f9", x"fc", x"fd", x"01", x"fd",
    x"fe", x"fd", x"fe", x"fc", x"02", x"02", x"ff", x"03",
    x"03", x"ff", x"fc", x"fc", x"ff", x"fe", x"fe", x"01",
    x"04", x"fb", x"fe", x"fd", x"ff", x"fc", x"fc", x"00",
    x"fb", x"fd", x"01", x"01", x"04", x"00", x"f9", x"02",
    x"03", x"04", x"03", x"fc", x"01", x"ff", x"fb", x"fc",
    x"fc", x"fe", x"01", x"02", x"01", x"ff", x"03", x"fc",
    x"00", x"fc", x"fb", x"fa", x"fb", x"fe", x"fc", x"fc",
    x"f6", x"fd", x"fe", x"fa", x"fe", x"fe", x"01", x"fb",
    x"04", x"fc", x"fe", x"fc", x"fe", x"f8", x"03", x"fc",
    x"f4", x"fc", x"f9", x"f9", x"ff", x"f9", x"00", x"fa",
    x"fa", x"00", x"f9", x"ff", x"fd", x"ff", x"fc", x"00",
    x"fd", x"f9", x"f6", x"fc", x"f9", x"00", x"fb", x"04",
    x"01", x"fb", x"fa", x"03", x"00", x"00", x"f5", x"fa",
    x"fc", x"04", x"fa", x"f9", x"fc", x"02", x"fd", x"f9",
    x"03", x"fc", x"01", x"00", x"fa", x"ff", x"fb", x"fb",
    x"02", x"03", x"fc", x"02", x"04", x"fd", x"fe", x"fb",
    x"04", x"03", x"ff", x"03", x"fc", x"fe", x"ff", x"ff",
    x"03", x"fa", x"02", x"00", x"00", x"01", x"fe", x"fa",
    x"fa", x"00", x"f9", x"f8", x"f8", x"fe", x"03", x"ff",
    x"f8", x"fe", x"fd", x"fb", x"fc", x"01", x"fb", x"fd",
    x"ff", x"fd", x"fd", x"fb", x"02", x"f6", x"00", x"00",
    x"fb", x"fc", x"00", x"fb", x"fd", x"01", x"ff", x"fc",
    x"02", x"fe", x"fb", x"02", x"fa", x"fb", x"fb", x"fc",
    x"fd", x"fd", x"00", x"03", x"03", x"fd", x"06", x"01",
    x"f7", x"ff", x"02", x"fc", x"fc", x"f8", x"06", x"03",
    x"fe", x"f6", x"fc", x"03", x"03", x"fc", x"04", x"f6",
    x"fc", x"f8", x"fa", x"fd", x"05", x"05", x"01", x"00",
    x"03", x"fd", x"04", x"00", x"fc", x"ff", x"01", x"03",
    x"fd", x"01", x"fd", x"fc", x"ff", x"01", x"01", x"fd",
    x"04", x"fc", x"fc", x"fb", x"01", x"fc", x"00", x"fc",
    x"05", x"00", x"04", x"02", x"04", x"02", x"fd", x"fd",
    x"fc", x"04", x"ff", x"01", x"f9", x"fa", x"fe", x"00",
    x"f9", x"ff", x"05", x"ff", x"fd", x"01", x"f6", x"f8",
    x"05", x"01", x"f8", x"00", x"01", x"f5", x"fb", x"fd",
    x"fa", x"00", x"fc", x"00", x"01", x"fb", x"f9", x"ff",
    x"ff", x"fd", x"fa", x"ff", x"ff", x"02", x"f8", x"fb",
    x"fa", x"fc", x"fc", x"fa", x"fe", x"01", x"ff", x"01",
    x"02", x"fe", x"00", x"fb", x"fc", x"fb", x"fd", x"fc",
    x"04", x"ff", x"01", x"fe", x"01", x"fe", x"00", x"ff",
    x"f9", x"04", x"ff", x"fc", x"fc", x"02", x"fb", x"fd",
    x"ff", x"01", x"f8", x"02", x"f5", x"fa", x"fc", x"ff",
    x"fe", x"02", x"fb", x"02", x"fc", x"fa", x"03", x"fe",
    x"01", x"03", x"00", x"fd", x"fc", x"01", x"04", x"01",
    x"fd", x"04", x"04", x"04", x"fe", x"ff", x"ff", x"fe",
    x"fd", x"fb", x"f9", x"fb", x"00", x"fb", x"04", x"fc",
    x"fb", x"04", x"fd", x"fd", x"01", x"00", x"ff", x"fc",
    x"fc", x"01", x"fd", x"fe", x"fa", x"fb", x"fd", x"fc",
    x"ff", x"fc", x"fe", x"00", x"01", x"f7", x"04", x"fd",
    x"04", x"fc", x"02", x"fd", x"fe", x"fd", x"f9", x"04",
    x"fe", x"ff", x"ff", x"01", x"fc", x"fc", x"f9", x"fa",
    x"03", x"ff", x"fe", x"04", x"fd", x"04", x"fd", x"ff",
    x"03", x"fd", x"00", x"01", x"ff", x"01", x"03", x"04",
    x"05", x"fd", x"fb", x"fd", x"fc", x"fb", x"fc", x"fc",
    x"fc", x"fe", x"ff", x"fd", x"fa", x"fe", x"00", x"fc",
    x"fc", x"ff", x"fa", x"04", x"00", x"fb", x"02", x"fe",
    x"01", x"ff", x"01", x"f8", x"fd", x"03", x"ff", x"fe",
    x"ff", x"f9", x"f6", x"fd", x"fd", x"fa", x"02", x"00",
    x"fc", x"04", x"01", x"01", x"00", x"fc", x"00", x"01",
    x"fd", x"ff", x"fe", x"fc", x"fe", x"fe", x"03", x"f7",
    x"fb", x"02", x"f8", x"04", x"fb", x"fd", x"03", x"00",
    x"fb", x"03", x"ff", x"fd", x"03", x"f7", x"fb", x"ff",
    x"04", x"f9", x"00", x"fe", x"fc", x"fa", x"02", x"fc",
    x"00", x"fe", x"01", x"02", x"04", x"00", x"ff", x"ff",
    x"f4", x"fd", x"fa", x"ff", x"ff", x"00", x"04", x"03",
    x"03", x"02", x"fc", x"fe", x"fe", x"01", x"fa", x"f8",
    x"02", x"01", x"fe", x"fa", x"f8", x"f6", x"fe", x"fb",
    x"fe", x"04", x"fd", x"ff", x"ff", x"00", x"ff", x"ff",
    x"02", x"fd", x"fc", x"fc", x"fc", x"01", x"fb", x"ff",
    x"ec", x"e1", x"14", x"07", x"19", x"e4", x"0d", x"f9",
    x"ae", x"78", x"2b", x"26", x"45", x"20", x"03", x"d5",
    x"fb", x"11", x"f2", x"df", x"c8", x"fa", x"02", x"07",
    x"07", x"20", x"2f", x"ee", x"e8", x"c2", x"e9", x"d0",
    x"cc", x"ec", x"d6", x"1d", x"02", x"df", x"04", x"15",
    x"2e", x"14", x"5d", x"1c", x"36", x"d4", x"15", x"29",
    x"f5", x"1e", x"18", x"f9", x"0d", x"24", x"4b", x"f5",
    x"05", x"e7", x"ea", x"0a", x"af", x"c1", x"bd", x"fe",
    x"35", x"26", x"46", x"3d", x"53", x"3c", x"3d", x"52",
    x"11", x"0d", x"0a", x"2f", x"f8", x"20", x"33", x"14",
    x"02", x"ed", x"fa", x"da", x"d7", x"c4", x"d2", x"a4",
    x"a5", x"d9", x"0e", x"00", x"12", x"19", x"09", x"16",
    x"72", x"f4", x"e8", x"0a", x"ee", x"f2", x"d5", x"f0",
    x"ed", x"a7", x"bf", x"a9", x"fe", x"09", x"5c", x"4a",
    x"2a", x"49", x"33", x"28", x"3b", x"e5", x"f2", x"0a",
    x"fa", x"0a", x"01", x"ee", x"f6", x"d7", x"e0", x"fa",
    x"dd", x"06", x"02", x"fc", x"ed", x"de", x"ea", x"e6",
    x"1c", x"5d", x"37", x"58", x"1b", x"45", x"44", x"22",
    x"2f", x"3c", x"2d", x"fb", x"fd", x"19", x"3a", x"02",
    x"eb", x"04", x"fc", x"03", x"fb", x"02", x"fc", x"03",
    x"fd", x"03", x"07", x"03", x"d0", x"d3", x"28", x"fd",
    x"16", x"3c", x"1f", x"f7", x"cc", x"e9", x"c0", x"cb",
    x"d1", x"bd", x"a6", x"fe", x"e9", x"ef", x"39", x"2c",
    x"3e", x"0c", x"25", x"33", x"e3", x"db", x"fa", x"13",
    x"e6", x"00", x"0b", x"34", x"49", x"3b", x"f1", x"ff",
    x"ca", x"f7", x"ee", x"0a", x"2e", x"14", x"e9", x"fe",
    x"00", x"27", x"d8", x"0c", x"28", x"34", x"1f", x"09",
    x"1a", x"c8", x"c1", x"2e", x"00", x"11", x"cd", x"f8",
    x"fa", x"00", x"12", x"31", x"05", x"20", x"19", x"c1",
    x"b6", x"fe", x"0d", x"fe", x"f4", x"2b", x"18", x"1d",
    x"74", x"0d", x"42", x"07", x"0a", x"01", x"ff", x"06",
    x"04", x"ff", x"07", x"01", x"18", x"d5", x"0c", x"1c",
    x"33", x"59", x"1d", x"50", x"1d", x"50", x"1c", x"e0",
    x"21", x"00", x"e8", x"14", x"f2", x"dc", x"f0", x"c9",
    x"dd", x"07", x"d0", x"ba", x"fb", x"d5", x"cb", x"18",
    x"2a", x"57", x"14", x"32", x"4b", x"57", x"37", x"16",
    x"01", x"01", x"f6", x"e8", x"00", x"11", x"de", x"f2",
    x"fa", x"d8", x"06", x"0f", x"0a", x"dc", x"e2", x"08",
    x"cb", x"da", x"0c", x"11", x"26", x"54", x"1c", x"2a",
    x"26", x"37", x"3f", x"f0", x"e2", x"16", x"f5", x"07",
    x"ee", x"e5", x"f7", x"c3", x"0e", x"01", x"fb", x"07",
    x"03", x"f8", x"00", x"04", x"01", x"3b", x"1d", x"31",
    x"4e", x"2f", x"0e", x"49", x"29", x"17", x"3a", x"b5",
    x"cb", x"20", x"e8", x"fe", x"ea", x"f8", x"fc", x"24",
    x"0a", x"ef", x"16", x"cb", x"8a", x"cf", x"ae", x"b4",
    x"fe", x"03", x"04", x"fd", x"05", x"fe", x"fb", x"fe",
    x"fd", x"e3", x"d6", x"bf", x"37", x"eb", x"da", x"0d",
    x"f8", x"e7", x"f5", x"e1", x"f1", x"0b", x"e1", x"d6",
    x"3e", x"f1", x"c6", x"28", x"e7", x"ef", x"27", x"d8",
    x"c5", x"28", x"cf", x"c4", x"33", x"fc", x"42", x"12",
    x"26", x"23", x"0a", x"11", x"31", x"48", x"08", x"36",
    x"1b", x"37", x"25", x"0d", x"0f", x"ec", x"fa", x"f1",
    x"fc", x"d8", x"ff", x"23", x"05", x"05", x"f9", x"0e",
    x"06", x"16", x"c3", x"eb", x"0a", x"07", x"ee", x"01",
    x"fa", x"fb", x"ff", x"fc", x"ff", x"ff", x"02", x"ff",
    x"ff", x"fb", x"f5", x"f9", x"fc", x"01", x"fc", x"fd",
    x"fc", x"00", x"4a", x"f9", x"08", x"12", x"3c", x"2e",
    x"1e", x"17", x"18", x"c1", x"cc", x"29", x"b4", x"bd",
    x"ed", x"dd", x"d2", x"d5", x"d4", x"12", x"04", x"07",
    x"07", x"ea", x"21", x"14", x"0b", x"e0", x"cf", x"04",
    x"e7", x"de", x"31", x"4b", x"84", x"3b", x"17", x"dc",
    x"14", x"d0", x"c5", x"ee", x"e7", x"ef", x"1c", x"1b",
    x"dd", x"c3", x"4a", x"f2", x"dd", x"dc", x"e5", x"e3",
    x"c8", x"db", x"eb", x"cb", x"fb", x"02", x"1c", x"4f",
    x"18", x"d0", x"f2", x"11", x"e7", x"d9", x"f4", x"c2",
    x"13", x"29", x"fa", x"a7", x"e3", x"15", x"4d", x"29",
    x"1d", x"4c", x"16", x"c4", x"19", x"18", x"06", x"0b",
    x"1a", x"49", x"14", x"3a", x"3d", x"13", x"e5", x"0a",
    x"e4", x"f0", x"2c", x"fa", x"cd", x"17", x"22", x"f1",
    x"0f", x"08", x"fc", x"ec", x"cf", x"ff", x"42", x"d8",
    x"b2", x"2d", x"09", x"e5", x"29", x"31", x"2c", x"3b",
    x"5a", x"34", x"26", x"04", x"2f", x"2e", x"12", x"42",
    x"f3", x"19", x"43", x"41", x"71", x"28", x"44", x"1c",
    x"79", x"23", x"28", x"28", x"2d", x"22", x"19", x"32",
    x"21", x"d7", x"73", x"50", x"29", x"11", x"21", x"fc",
    x"d3", x"ba", x"a4", x"d8", x"d2", x"f8", x"f3", x"dc",
    x"1d", x"de", x"c0", x"f1", x"19", x"1f", x"21", x"10",
    x"00", x"0d", x"fa", x"df", x"c1", x"4f", x"e1", x"ac",
    x"dc", x"e9", x"cc", x"0a", x"fb", x"b7", x"e4", x"12",
    x"02", x"f6", x"16", x"02", x"a7", x"a7", x"ed", x"9f",
    x"b6", x"0d", x"ef", x"03", x"e7", x"22", x"25", x"f0",
    x"de", x"d6", x"16", x"01", x"1c", x"3b", x"1d", x"2f",
    x"39", x"19", x"ee", x"d2", x"f2", x"fb", x"fa", x"d2",
    x"01", x"24", x"83", x"43", x"39", x"36", x"2e", x"2c",
    x"44", x"ca", x"ca", x"d6", x"1e", x"29", x"13", x"e4",
    x"ec", x"38", x"e8", x"bd", x"b9", x"ee", x"ea", x"20",
    x"35", x"1b", x"ff", x"07", x"14", x"45", x"63", x"8f",
    x"00", x"e5", x"1b", x"cd", x"ba", x"d8", x"38", x"06",
    x"0c", x"b9", x"dd", x"d6", x"a1", x"c7", x"e4", x"f2",
    x"04", x"00", x"ed", x"e4", x"fa", x"ba", x"e4", x"d8",
    x"ba", x"91", x"b6", x"fc", x"cd", x"d5", x"f1", x"11",
    x"14", x"ff", x"02", x"04", x"00", x"fb", x"fc", x"fa",
    x"01", x"fb", x"09", x"12", x"09", x"cc", x"bf", x"d8",
    x"13", x"15", x"14", x"39", x"17", x"14", x"f1", x"d4",
    x"e0", x"eb", x"f7", x"36", x"2f", x"6a", x"57", x"25",
    x"f4", x"de", x"17", x"0c", x"f9", x"ef", x"f0", x"0b",
    x"16", x"18", x"39", x"17", x"04", x"c1", x"ec", x"06",
    x"f3", x"f1", x"f0", x"f0", x"37", x"58", x"0a", x"1e",
    x"f3", x"02", x"23", x"00", x"03", x"44", x"14", x"0a",
    x"2a", x"33", x"3e", x"77", x"15", x"e3", x"87", x"05",
    x"fc", x"1f", x"ea", x"e2", x"27", x"0e", x"fb", x"1d",
    x"f3", x"d2", x"18", x"f5", x"e8", x"0d", x"11", x"2d",
    x"22", x"2d", x"d6", x"02", x"05", x"fb", x"ff", x"fd",
    x"04", x"fe", x"fb", x"04", x"18", x"f0", x"eb", x"e5",
    x"f4", x"16", x"f1", x"de", x"fc", x"0b", x"ea", x"1c",
    x"21", x"1c", x"11", x"0b", x"f5", x"39", x"0a", x"eb",
    x"2c", x"9f", x"da", x"e4", x"59", x"bf", x"00", x"eb",
    x"d6", x"ea", x"e8", x"01", x"0e", x"04", x"0f", x"12",
    x"e1", x"fa", x"3c", x"05", x"d2", x"e9", x"0a", x"e5",
    x"9a", x"05", x"bf", x"99", x"fe", x"f6", x"fd", x"f8",
    x"34", x"1b", x"fe", x"12", x"06", x"f4", x"e1", x"0a",
    x"f0", x"01", x"c6", x"b1", x"fa", x"f3", x"2f", x"14",
    x"19", x"54", x"0f", x"1b", x"fe", x"08", x"08", x"fe",
    x"0c", x"0c", x"03", x"0c", x"08", x"20", x"03", x"14",
    x"10", x"f4", x"d3", x"04", x"f3", x"b9", x"53", x"14",
    x"05", x"58", x"fc", x"15", x"63", x"ef", x"0d", x"0f",
    x"13", x"ec", x"ff", x"fb", x"08", x"13", x"e7", x"fc",
    x"fc", x"fe", x"04", x"01", x"01", x"fe", x"05", x"08",
    x"fe", x"2d", x"0e", x"39", x"e5", x"f9", x"ff", x"ef",
    x"f0", x"fb", x"ae", x"ed", x"13", x"e9", x"22", x"31",
    x"18", x"0a", x"fe", x"43", x"13", x"0e", x"1c", x"0c",
    x"05", x"2f", x"f5", x"17", x"22", x"38", x"2f", x"cc",
    x"49", x"47", x"ef", x"e1", x"ee", x"07", x"f7", x"22",
    x"d4", x"03", x"37", x"1a", x"44", x"6e", x"8d", x"42",
    x"36", x"01", x"e4", x"fc", x"d7", x"01", x"37", x"3d",
    x"03", x"07", x"2e", x"e2", x"06", x"df", x"f6", x"eb",
    x"02", x"fd", x"03", x"fe", x"fc", x"fd", x"fa", x"fb",
    x"fa", x"02", x"f9", x"fd", x"ff", x"01", x"02", x"02",
    x"fe", x"fe", x"35", x"ee", x"e0", x"40", x"2a", x"45",
    x"35", x"1a", x"d9", x"23", x"f8", x"21", x"fc", x"bc",
    x"7b", x"07", x"a4", x"96", x"6a", x"5a", x"1a", x"e6",
    x"db", x"ef", x"25", x"f5", x"27", x"d5", x"06", x"06",
    x"12", x"0f", x"0f", x"48", x"09", x"c6", x"f7", x"12",
    x"f9", x"ed", x"21", x"0c", x"ef", x"08", x"00", x"20",
    x"42", x"41", x"20", x"f2", x"c2", x"b2", x"c3", x"02",
    x"18", x"25", x"39", x"2e", x"04", x"ea", x"c3", x"de",
    x"07", x"11", x"05", x"13", x"4a", x"3b", x"27", x"e3",
    x"1d", x"e8", x"04", x"0f", x"0a", x"f4", x"11", x"f4",
    x"f4", x"f3", x"ed", x"23", x"16", x"fb", x"08", x"01",
    x"fc", x"f4", x"e4", x"e6", x"00", x"d9", x"a1", x"14",
    x"26", x"1d", x"11", x"18", x"03", x"02", x"09", x"28",
    x"f2", x"16", x"20", x"1c", x"20", x"11", x"a7", x"f7",
    x"10", x"12", x"21", x"03", x"4c", x"27", x"e6", x"1a",
    x"f3", x"0a", x"01", x"f8", x"f9", x"1e", x"22", x"ea",
    x"b9", x"c2", x"69", x"18", x"09", x"b6", x"c9", x"f3",
    x"24", x"f7", x"2d", x"20", x"02", x"1d", x"19", x"c4",
    x"e3", x"de", x"a8", x"df", x"8d", x"e3", x"dc", x"c6",
    x"2d", x"3c", x"42", x"05", x"0d", x"36", x"16", x"0a",
    x"0e", x"cf", x"bb", x"b1", x"d7", x"ff", x"05", x"c0",
    x"d6", x"eb", x"16", x"fa", x"2b", x"1f", x"28", x"bc",
    x"03", x"fa", x"c7", x"d0", x"fb", x"47", x"f2", x"01",
    x"06", x"ef", x"fb", x"e5", x"bd", x"ea", x"f3", x"46",
    x"ff", x"e5", x"f7", x"41", x"03", x"c8", x"dc", x"26",
    x"f1", x"c2", x"7b", x"07", x"47", x"2d", x"f3", x"f0",
    x"06", x"06", x"3b", x"25", x"33", x"31", x"2b", x"0b",
    x"f4", x"01", x"ea", x"14", x"04", x"57", x"e0", x"fa",
    x"44", x"0e", x"ba", x"13", x"c7", x"dc", x"49", x"45",
    x"2c", x"d2", x"23", x"16", x"ce", x"aa", x"bd", x"b2",
    x"e1", x"34", x"69", x"ad", x"e1", x"e2", x"95", x"9a",
    x"fc", x"15", x"26", x"0b", x"02", x"26", x"f8", x"d1",
    x"ef", x"12", x"f7", x"ee", x"e1", x"fe", x"f3", x"ed",
    x"16", x"f6", x"31", x"27", x"28", x"16", x"2f", x"2e",
    x"1b", x"df", x"95", x"f1", x"01", x"e6", x"0b", x"01",
    x"eb", x"fe", x"03", x"fc", x"02", x"01", x"04", x"fd",
    x"04", x"05", x"d2", x"c7", x"c4", x"28", x"e5", x"ba",
    x"41", x"28", x"14", x"0a", x"c6", x"da", x"f9", x"fd",
    x"19", x"16", x"22", x"ec", x"ff", x"24", x"ff", x"2f",
    x"2b", x"2f", x"fb", x"cd", x"ba", x"ed", x"c0", x"cb",
    x"e7", x"10", x"14", x"5d", x"47", x"0e", x"f3", x"cb",
    x"a1", x"08", x"d6", x"be", x"2d", x"32", x"2d", x"f3",
    x"0d", x"f8", x"01", x"f7", x"f2", x"1d", x"32", x"59",
    x"44", x"9d", x"3e", x"4f", x"e3", x"ee", x"f5", x"0c",
    x"30", x"fc", x"ff", x"d6", x"3a", x"29", x"19", x"2b",
    x"f7", x"8f", x"df", x"d1", x"a1", x"f8", x"ee", x"07",
    x"3b", x"5f", x"3d", x"fc", x"02", x"fc", x"03", x"05",
    x"01", x"fe", x"03", x"00", x"b9", x"ba", x"2c", x"0a",
    x"00", x"19", x"3c", x"23", x"11", x"17", x"23", x"89",
    x"a5", x"d3", x"22", x"30", x"37", x"14", x"ac", x"dc",
    x"9b", x"f7", x"eb", x"13", x"e7", x"dd", x"97", x"c2",
    x"ce", x"ba", x"d3", x"f7", x"20", x"e9", x"d7", x"09",
    x"f4", x"fe", x"f4", x"db", x"cd", x"e1", x"19", x"07",
    x"eb", x"0e", x"02", x"df", x"28", x"04", x"06", x"09",
    x"d8", x"fd", x"c8", x"d0", x"0c", x"5d", x"12", x"f6",
    x"07", x"1f", x"22", x"d1", x"a8", x"cc", x"17", x"cc",
    x"20", x"cd", x"29", x"2a", x"fb", x"05", x"fe", x"0c",
    x"08", x"04", x"0d", x"00", x"05", x"e9", x"ec", x"e9",
    x"54", x"30", x"03", x"17", x"10", x"fa", x"07", x"a0",
    x"9d", x"f2", x"b1", x"b0", x"33", x"2f", x"18", x"4b",
    x"2c", x"04", x"56", x"d8", x"dd", x"fa", x"dc", x"ec",
    x"05", x"fe", x"04", x"02", x"01", x"00", x"02", x"02",
    x"02", x"d6", x"c6", x"6e", x"e0", x"e8", x"cd", x"fe",
    x"19", x"20", x"e3", x"a3", x"8b", x"03", x"f4", x"ff",
    x"f7", x"e6", x"df", x"c7", x"bf", x"b4", x"22", x"ff",
    x"0c", x"4e", x"e3", x"d7", x"a4", x"34", x"ef", x"fa",
    x"11", x"31", x"02", x"37", x"46", x"7c", x"51", x"92",
    x"ab", x"18", x"0a", x"c8", x"fc", x"f7", x"0a", x"e2",
    x"ca", x"07", x"e8", x"c6", x"02", x"22", x"44", x"02",
    x"ea", x"e5", x"e3", x"28", x"20", x"55", x"2d", x"08",
    x"02", x"fc", x"01", x"fc", x"fd", x"fc", x"01", x"05",
    x"fb", x"fe", x"fe", x"03", x"fd", x"01", x"01", x"01",
    x"ff", x"03", x"e5", x"f2", x"cc", x"53", x"3f", x"18",
    x"ee", x"0f", x"23", x"f8", x"c7", x"f8", x"0f", x"f3",
    x"e5", x"05", x"eb", x"1c", x"1c", x"fa", x"cb", x"09",
    x"01", x"15", x"25", x"20", x"25", x"e5", x"df", x"cf",
    x"f3", x"e0", x"26", x"05", x"02", x"1e", x"ee", x"d6",
    x"e8", x"39", x"35", x"17", x"34", x"1f", x"00", x"32",
    x"c8", x"bb", x"41", x"05", x"07", x"ac", x"fb", x"13",
    x"03", x"cf", x"f4", x"3a", x"df", x"d6", x"9f", x"a6",
    x"b4", x"10", x"00", x"f8", x"0a", x"27", x"18", x"b3",
    x"bc", x"bc", x"ad", x"94", x"9f", x"17", x"1e", x"0d",
    x"f4", x"f5", x"0f", x"bc", x"d7", x"f8", x"0a", x"f8",
    x"f8", x"0d", x"17", x"1a", x"0d", x"03", x"8a", x"35",
    x"0a", x"f4", x"28", x"06", x"f4", x"2f", x"37", x"fb",
    x"0b", x"f7", x"11", x"fe", x"ad", x"d1", x"01", x"9e",
    x"89", x"cc", x"8a", x"b8", x"ae", x"ef", x"f5", x"c9",
    x"af", x"e2", x"f2", x"f0", x"06", x"c5", x"15", x"04",
    x"f4", x"e1", x"e7", x"ef", x"ca", x"e1", x"f8", x"15",
    x"3a", x"05", x"dc", x"03", x"fe", x"03", x"04", x"23",
    x"bd", x"9d", x"ea", x"db", x"b4", x"d5", x"24", x"fd",
    x"02", x"10", x"10", x"00", x"22", x"15", x"11", x"29",
    x"46", x"df", x"f7", x"12", x"ff", x"e5", x"ee", x"ed",
    x"db", x"c0", x"fa", x"fe", x"f5", x"e4", x"17", x"40",
    x"07", x"e8", x"df", x"21", x"dc", x"40", x"fa", x"e6",
    x"e6", x"2a", x"02", x"fb", x"59", x"24", x"19", x"1a",
    x"35", x"21", x"02", x"0c", x"e0", x"eb", x"00", x"1a",
    x"17", x"19", x"0c", x"f9", x"e6", x"e0", x"e6", x"e4",
    x"d2", x"f5", x"eb", x"fd", x"18", x"21", x"18", x"fb",
    x"05", x"ee", x"fa", x"d9", x"dc", x"55", x"19", x"10",
    x"07", x"0b", x"d3", x"36", x"dc", x"d8", x"12", x"11",
    x"28", x"07", x"12", x"3b", x"08", x"1a", x"1b", x"ea",
    x"bf", x"87", x"29", x"fa", x"e8", x"da", x"d1", x"f6",
    x"f5", x"0a", x"22", x"f7", x"f3", x"ff", x"ec", x"e8",
    x"ef", x"23", x"06", x"0d", x"e0", x"eb", x"02", x"ec",
    x"ce", x"a4", x"e9", x"e0", x"f6", x"f6", x"db", x"f6",
    x"29", x"0e", x"1a", x"e6", x"e5", x"f6", x"f4", x"1c",
    x"02", x"04", x"ff", x"ff", x"ff", x"03", x"00", x"fb",
    x"fb", x"fb", x"e8", x"f0", x"ef", x"ad", x"f1", x"e9",
    x"29", x"11", x"0c", x"b7", x"dd", x"ff", x"f8", x"14",
    x"16", x"2c", x"1f", x"49", x"e3", x"eb", x"19", x"f0",
    x"0d", x"1c", x"fa", x"00", x"e9", x"d5", x"e7", x"e0",
    x"1e", x"0d", x"f0", x"3a", x"16", x"1b", x"03", x"06",
    x"03", x"fa", x"e6", x"f3", x"18", x"0c", x"14", x"df",
    x"de", x"fc", x"f7", x"dd", x"d4", x"15", x"e6", x"e1",
    x"32", x"b8", x"cc", x"28", x"c4", x"01", x"0a", x"db",
    x"de", x"e2", x"d2", x"e7", x"17", x"02", x"0b", x"13",
    x"fa", x"d9", x"d3", x"e5", x"cf", x"0d", x"f3", x"08",
    x"0c", x"02", x"48", x"fe", x"03", x"ff", x"00", x"fc",
    x"ff", x"05", x"02", x"fb", x"3a", x"e4", x"0b", x"34",
    x"18", x"e9", x"00", x"15", x"fd", x"33", x"d6", x"f2",
    x"06", x"12", x"0f", x"4d", x"32", x"03", x"eb", x"f7",
    x"ed", x"df", x"0c", x"fa", x"f9", x"c5", x"bc", x"0b",
    x"27", x"10", x"d8", x"ca", x"e9", x"ee", x"05", x"19",
    x"03", x"f7", x"e5", x"10", x"f8", x"cc", x"b7", x"f9",
    x"11", x"0d", x"f3", x"00", x"21", x"15", x"03", x"ed",
    x"f5", x"16", x"1a", x"ff", x"07", x"62", x"eb", x"e2",
    x"ee", x"25", x"14", x"17", x"11", x"c1", x"1e", x"21",
    x"1e", x"1c", x"03", x"1f", x"01", x"01", x"fa", x"f9",
    x"fe", x"fe", x"07", x"02", x"f8", x"0c", x"05", x"02",
    x"09", x"11", x"1f", x"0e", x"1f", x"19", x"0d", x"26",
    x"09", x"2d", x"d7", x"ec", x"13", x"f6", x"dd", x"1b",
    x"fe", x"e9", x"04", x"e3", x"fb", x"18", x"0c", x"0a",
    x"02", x"fb", x"03", x"04", x"03", x"fc", x"02", x"fb",
    x"fc", x"e9", x"c8", x"a5", x"0f", x"07", x"1c", x"09",
    x"01", x"03", x"fb", x"37", x"0e", x"db", x"ac", x"dc",
    x"f0", x"fe", x"dd", x"ec", x"dc", x"ec", x"00", x"10",
    x"05", x"0a", x"fd", x"e6", x"c9", x"f2", x"05", x"f9",
    x"1f", x"4b", x"30", x"3e", x"25", x"27", x"07", x"02",
    x"ca", x"c4", x"f4", x"d2", x"e8", x"02", x"d5", x"e2",
    x"41", x"dc", x"da", x"f1", x"13", x"ea", x"f4", x"da",
    x"ef", x"1d", x"10", x"07", x"19", x"33", x"0f", x"08",
    x"fc", x"fe", x"ff", x"05", x"04", x"fb", x"04", x"fd",
    x"fe", x"fa", x"fe", x"02", x"fb", x"fc", x"01", x"ff",
    x"02", x"fc", x"53", x"45", x"17", x"e9", x"a5", x"d7",
    x"ca", x"d1", x"e0", x"14", x"f5", x"3d", x"de", x"08",
    x"e7", x"f0", x"ee", x"fc", x"c4", x"e2", x"22", x"19",
    x"3e", x"2c", x"10", x"1d", x"17", x"0d", x"d7", x"ea",
    x"06", x"fb", x"f0", x"0e", x"05", x"2a", x"34", x"b9",
    x"d4", x"2b", x"13", x"ea", x"0c", x"0d", x"04", x"0f",
    x"d2", x"dd", x"17", x"f7", x"f9", x"14", x"3c", x"0e",
    x"0f", x"ec", x"00", x"f9", x"0a", x"03", x"06", x"fe",
    x"f5", x"2b", x"d5", x"f3", x"e3", x"03", x"1a", x"e6",
    x"e5", x"b9", x"ec", x"ea", x"d7", x"09", x"e3", x"08",
    x"19", x"24", x"1e", x"fe", x"1a", x"fd", x"0d", x"fd",
    x"09", x"1d", x"04", x"1b", x"1c", x"3f", x"32", x"16",
    x"ed", x"10", x"0f", x"2f", x"21", x"c9", x"f7", x"08",
    x"0a", x"f6", x"0c", x"22", x"38", x"f4", x"36", x"ed",
    x"19", x"22", x"d5", x"b7", x"e3", x"c1", x"c6", x"02",
    x"04", x"26", x"cf", x"28", x"67", x"ef", x"2c", x"1b",
    x"01", x"07", x"3c", x"24", x"1f", x"b2", x"3b", x"f2",
    x"cb", x"1a", x"0a", x"ec", x"4d", x"31", x"22", x"3e",
    x"b2", x"7f", x"0f", x"19", x"12", x"03", x"e8", x"97",
    x"e1", x"af", x"a6", x"9e", x"65", x"a9", x"e1", x"09",
    x"04", x"ef", x"08", x"eb", x"1b", x"25", x"07", x"fe",
    x"33", x"39", x"1e", x"0c", x"c3", x"fd", x"f6", x"26",
    x"e8", x"bb", x"77", x"2d", x"9c", x"9b", x"0e", x"2e",
    x"f3", x"04", x"00", x"e7", x"f0", x"fc", x"23", x"c4",
    x"b9", x"64", x"df", x"e7", x"2e", x"1d", x"2a", x"56",
    x"c9", x"ca", x"fe", x"ea", x"f1", x"3f", x"22", x"00",
    x"46", x"d5", x"e7", x"f0", x"c9", x"0b", x"23", x"d7",
    x"f6", x"29", x"09", x"cc", x"d6", x"b9", x"d9", x"ef",
    x"04", x"e1", x"0c", x"ff", x"f1", x"f2", x"dc", x"d8",
    x"b5", x"01", x"04", x"ce", x"e4", x"fa", x"05", x"5c",
    x"17", x"22", x"fd", x"f2", x"07", x"17", x"40", x"31",
    x"16", x"00", x"24", x"f6", x"e6", x"40", x"2f", x"19",
    x"18", x"2c", x"3c", x"f2", x"23", x"20", x"38", x"ec",
    x"0b", x"f4", x"e8", x"41", x"0b", x"08", x"21", x"24",
    x"e7", x"ec", x"f6", x"f3", x"ed", x"05", x"d1", x"d4",
    x"0e", x"03", x"00", x"fe", x"03", x"fe", x"00", x"02",
    x"fd", x"02", x"29", x"f0", x"3f", x"e4", x"eb", x"ea",
    x"0e", x"f8", x"fd", x"02", x"fb", x"13", x"dd", x"c3",
    x"d5", x"ef", x"24", x"49", x"16", x"28", x"0b", x"17",
    x"06", x"17", x"ff", x"f8", x"33", x"ef", x"d7", x"c9",
    x"c6", x"e5", x"16", x"dd", x"09", x"e3", x"e3", x"d5",
    x"f9", x"d6", x"cf", x"00", x"94", x"8e", x"f9", x"2a",
    x"13", x"0f", x"f5", x"12", x"fe", x"ed", x"e8", x"da",
    x"37", x"4f", x"3c", x"36", x"2f", x"0c", x"4c", x"a4",
    x"e2", x"24", x"fb", x"e4", x"45", x"28", x"22", x"42",
    x"24", x"aa", x"19", x"0e", x"1c", x"fc", x"ee", x"03",
    x"ed", x"d0", x"92", x"06", x"fb", x"fb", x"0b", x"ff",
    x"09", x"02", x"fd", x"06", x"c7", x"f3", x"24", x"e2",
    x"e7", x"0a", x"dd", x"16", x"3b", x"27", x"f4", x"1f",
    x"2a", x"1c", x"db", x"06", x"2a", x"10", x"f2", x"07",
    x"06", x"f3", x"01", x"f8", x"ca", x"07", x"bc", x"d9",
    x"d4", x"e0", x"09", x"ec", x"07", x"20", x"20", x"49",
    x"30", x"1a", x"1c", x"3a", x"02", x"d3", x"08", x"c6",
    x"8c", x"f0", x"e0", x"e8", x"f6", x"e8", x"0f", x"1d",
    x"34", x"54", x"15", x"0b", x"14", x"20", x"33", x"fc",
    x"43", x"41", x"d1", x"f1", x"e0", x"b9", x"05", x"1c",
    x"48", x"ef", x"71", x"47", x"fc", x"f0", x"fd", x"fc",
    x"fc", x"f4", x"f5", x"f0", x"f5", x"f4", x"18", x"e5",
    x"20", x"13", x"12", x"00", x"36", x"00", x"35", x"c7",
    x"d7", x"47", x"b6", x"ef", x"ec", x"c4", x"df", x"1f",
    x"0f", x"05", x"f6", x"cf", x"cd", x"12", x"bb", x"a1",
    x"01", x"fc", x"ff", x"03", x"fd", x"fc", x"fe", x"fe",
    x"00", x"1a", x"02", x"19", x"18", x"f7", x"13", x"fb",
    x"37", x"1f", x"00", x"12", x"e1", x"f3", x"f4", x"24",
    x"10", x"0a", x"1c", x"f5", x"dc", x"e3", x"03", x"38",
    x"4c", x"11", x"60", x"1b", x"dd", x"d2", x"e1", x"ef",
    x"12", x"1a", x"05", x"ff", x"e1", x"fc", x"1d", x"50",
    x"eb", x"f3", x"fa", x"ea", x"c9", x"f4", x"31", x"69",
    x"3d", x"1c", x"f6", x"aa", x"d0", x"04", x"03", x"40",
    x"20", x"f1", x"23", x"fe", x"b2", x"f5", x"e1", x"d0",
    x"fe", x"fa", x"00", x"f8", x"00", x"ff", x"fa", x"fa",
    x"f7", x"03", x"05", x"00", x"fd", x"00", x"fe", x"fb",
    x"fe", x"01", x"16", x"2a", x"23", x"1e", x"25", x"25",
    x"0b", x"fd", x"f4", x"2e", x"29", x"bb", x"22", x"e0",
    x"e4", x"f4", x"d6", x"fc", x"13", x"f8", x"12", x"08",
    x"00", x"e9", x"05", x"18", x"00", x"0f", x"1b", x"28",
    x"1a", x"08", x"02", x"f9", x"ee", x"1e", x"ec", x"e3",
    x"e6", x"f5", x"b4", x"dd", x"cd", x"e8", x"da", x"54",
    x"4c", x"35", x"35", x"e6", x"c4", x"1e", x"ee", x"fc",
    x"22", x"09", x"e6", x"3c", x"99", x"e4", x"2a", x"ac",
    x"ed", x"19", x"30", x"22", x"3f", x"14", x"07", x"2b",
    x"51", x"b6", x"dc", x"09", x"1a", x"f5", x"dd", x"ca",
    x"34", x"03", x"f8", x"0b", x"f4", x"02", x"1f", x"ea",
    x"ed", x"0e", x"fa", x"d0", x"07", x"2d", x"55", x"ea",
    x"4f", x"3f", x"df", x"12", x"2b", x"db", x"eb", x"10",
    x"cc", x"41", x"3b", x"ea", x"4e", x"1e", x"12", x"53",
    x"71", x"0f", x"28", x"35", x"0a", x"d0", x"c9", x"10",
    x"23", x"31", x"16", x"fc", x"0c", x"54", x"e4", x"01",
    x"ff", x"01", x"fe", x"01", x"f8", x"00", x"fe", x"02",
    x"fc", x"03", x"fc", x"fd", x"fa", x"fd", x"f8", x"fe",
    x"00", x"fd", x"fb", x"fc", x"02", x"fd", x"fd", x"ff",
    x"01", x"fa", x"01", x"f8", x"fc", x"fc", x"00", x"f9",
    x"fb", x"f8", x"00", x"f9", x"fd", x"fa", x"fa", x"fa",
    x"fb", x"00", x"f9", x"ff", x"fd", x"00", x"ff", x"fe",
    x"f9", x"f6", x"00", x"fd", x"01", x"02", x"02", x"fc",
    x"f7", x"00", x"05", x"f9", x"01", x"fb", x"03", x"03",
    x"fc", x"01", x"fe", x"00", x"02", x"fa", x"fc", x"04",
    x"fd", x"fd", x"fc", x"fb", x"03", x"01", x"ff", x"fc",
    x"03", x"05", x"fc", x"02", x"f9", x"fc", x"01", x"ff",
    x"fc", x"03", x"02", x"03", x"ff", x"fc", x"fa", x"ff",
    x"01", x"00", x"fa", x"04", x"fa", x"fe", x"fc", x"06",
    x"04", x"02", x"04", x"fa", x"02", x"02", x"ff", x"04",
    x"ff", x"fe", x"02", x"03", x"00", x"fb", x"fa", x"ff",
    x"fc", x"f6", x"ff", x"fe", x"fc", x"01", x"fd", x"ff",
    x"fd", x"fd", x"01", x"03", x"03", x"fb", x"fc", x"fc",
    x"fd", x"00", x"fa", x"fc", x"02", x"fe", x"f6", x"fe",
    x"fb", x"02", x"fe", x"ff", x"01", x"fe", x"00", x"fe",
    x"fa", x"01", x"02", x"ff", x"00", x"00", x"05", x"fb",
    x"03", x"fe", x"fb", x"f7", x"ff", x"fd", x"fc", x"fe",
    x"fa", x"fd", x"00", x"ff", x"ff", x"fe", x"f8", x"f4",
    x"fe", x"ff", x"00", x"f7", x"f9", x"ff", x"fe", x"ff",
    x"fa", x"ff", x"09", x"fe", x"00", x"04", x"00", x"fb",
    x"fc", x"02", x"f8", x"04", x"00", x"03", x"02", x"03",
    x"fb", x"fd", x"fa", x"01", x"f9", x"ff", x"04", x"04",
    x"02", x"f9", x"fb", x"f8", x"01", x"fb", x"f9", x"fe",
    x"04", x"fd", x"ff", x"03", x"fb", x"02", x"0a", x"02",
    x"fb", x"03", x"ff", x"fc", x"04", x"fd", x"fd", x"04",
    x"04", x"02", x"ff", x"f9", x"fe", x"fc", x"f5", x"ff",
    x"02", x"00", x"ff", x"ff", x"fd", x"04", x"01", x"02",
    x"01", x"fd", x"02", x"01", x"fd", x"02", x"fc", x"fb",
    x"f9", x"fe", x"f9", x"fa", x"fe", x"03", x"00", x"fa",
    x"fd", x"00", x"fe", x"fe", x"fd", x"ff", x"fc", x"fc",
    x"f9", x"fc", x"fe", x"00", x"fd", x"fe", x"fc", x"03",
    x"fd", x"03", x"f8", x"00", x"fd", x"f9", x"fe", x"f9",
    x"fc", x"02", x"ff", x"ff", x"fb", x"00", x"fc", x"fa",
    x"01", x"f7", x"fe", x"f4", x"00", x"05", x"fe", x"02",
    x"f5", x"fd", x"02", x"fa", x"fd", x"03", x"ff", x"01",
    x"04", x"ff", x"fd", x"05", x"f5", x"fb", x"01", x"03",
    x"00", x"00", x"fd", x"03", x"fd", x"fe", x"fe", x"ff",
    x"fd", x"02", x"00", x"02", x"fe", x"fc", x"fb", x"fb",
    x"fb", x"fd", x"00", x"f9", x"ff", x"fb", x"00", x"fa",
    x"02", x"02", x"fc", x"02", x"fb", x"03", x"f8", x"01",
    x"fc", x"01", x"ff", x"00", x"fc", x"f8", x"fd", x"fd",
    x"02", x"fe", x"04", x"01", x"fb", x"03", x"00", x"fd",
    x"ff", x"02", x"fc", x"fc", x"fa", x"fe", x"00", x"fb",
    x"f7", x"fb", x"00", x"ff", x"fc", x"f9", x"00", x"01",
    x"02", x"fd", x"fd", x"01", x"ff", x"f9", x"00", x"02",
    x"01", x"fe", x"fd", x"01", x"fc", x"fb", x"fc", x"fb",
    x"00", x"fd", x"ff", x"fe", x"fb", x"fe", x"00", x"00",
    x"03", x"fa", x"fc", x"fe", x"f8", x"fe", x"fa", x"f8",
    x"00", x"f8", x"f8", x"fe", x"ff", x"fa", x"fc", x"fb",
    x"02", x"f8", x"f8", x"ff", x"fd", x"fc", x"fe", x"fc",
    x"fc", x"fe", x"fe", x"03", x"fd", x"fc", x"fd", x"02",
    x"05", x"fc", x"04", x"01", x"fb", x"01", x"fb", x"00",
    x"00", x"02", x"02", x"02", x"fc", x"fe", x"02", x"f8",
    x"02", x"00", x"fc", x"fe", x"fd", x"ff", x"fc", x"f9",
    x"04", x"f9", x"fe", x"fa", x"fc", x"f8", x"fc", x"fd",
    x"f9", x"fc", x"04", x"fd", x"fc", x"fe", x"fc", x"fe",
    x"fb", x"fe", x"ff", x"03", x"fc", x"fb", x"fa", x"fb",
    x"fb", x"fb", x"fc", x"fe", x"00", x"fe", x"fa", x"ff",
    x"fc", x"f7", x"f7", x"fb", x"f8", x"00", x"fb", x"fd",
    x"04", x"fe", x"fe", x"04", x"f9", x"00", x"01", x"fd",
    x"02", x"f6", x"fb", x"fa", x"fb", x"01", x"f7", x"01",
    x"f9", x"01", x"fb", x"02", x"fa", x"f8", x"fe", x"fe",
    x"03", x"fe", x"01", x"07", x"fc", x"ff", x"fb", x"f9",
    x"01", x"04", x"fe", x"fc", x"02", x"02", x"f9", x"01",
    x"00", x"00", x"fa", x"fa", x"00", x"00", x"fd", x"fc",
    x"fb", x"ff", x"fd", x"02", x"f5", x"fc", x"01", x"fa",
    x"fd", x"fc", x"fd", x"00", x"02", x"fe", x"fa", x"ff",
    x"00", x"03", x"f9", x"03", x"fa", x"ff", x"fa", x"fe",
    x"2f", x"f3", x"f5", x"1f", x"af", x"02", x"dc", x"e5",
    x"c9", x"06", x"06", x"f9", x"05", x"02", x"dc", x"0c",
    x"cd", x"94", x"67", x"8f", x"c4", x"c3", x"de", x"f1",
    x"f5", x"05", x"ef", x"c2", x"b4", x"ed", x"9c", x"ea",
    x"26", x"20", x"2a", x"1f", x"cf", x"b4", x"f2", x"b3",
    x"a6", x"bd", x"f0", x"cd", x"ce", x"aa", x"01", x"14",
    x"e9", x"f3", x"d3", x"30", x"1e", x"fb", x"41", x"11",
    x"b0", x"6a", x"18", x"3c", x"f7", x"13", x"1b", x"01",
    x"16", x"e6", x"2c", x"3e", x"41", x"19", x"06", x"ec",
    x"e8", x"15", x"eb", x"11", x"f4", x"ed", x"c3", x"9f",
    x"8f", x"10", x"19", x"15", x"e6", x"fa", x"fb", x"d7",
    x"fc", x"e1", x"25", x"04", x"ec", x"bf", x"f9", x"11",
    x"e4", x"fe", x"0e", x"33", x"ed", x"f5", x"33", x"f3",
    x"11", x"03", x"0e", x"11", x"39", x"14", x"ce", x"ff",
    x"cf", x"ca", x"fb", x"8e", x"c2", x"da", x"d7", x"b5",
    x"dc", x"06", x"3e", x"16", x"23", x"03", x"1e", x"03",
    x"08", x"db", x"11", x"0b", x"3a", x"25", x"38", x"64",
    x"ff", x"ee", x"a8", x"02", x"2e", x"01", x"ea", x"e3",
    x"23", x"26", x"49", x"29", x"0b", x"d1", x"c6", x"ad",
    x"da", x"fd", x"02", x"02", x"fa", x"fc", x"fe", x"05",
    x"01", x"fe", x"cf", x"f8", x"0d", x"ec", x"02", x"05",
    x"04", x"2c", x"f7", x"07", x"00", x"24", x"0c", x"30",
    x"10", x"3e", x"20", x"f0", x"d6", x"e3", x"05", x"17",
    x"fd", x"23", x"10", x"0d", x"0a", x"26", x"f8", x"d4",
    x"f7", x"02", x"09", x"95", x"89", x"c4", x"30", x"28",
    x"1b", x"19", x"da", x"c1", x"b4", x"d2", x"e8", x"f3",
    x"24", x"f6", x"02", x"f6", x"f9", x"c8", x"b0", x"d2",
    x"18", x"dd", x"e3", x"92", x"cf", x"0f", x"dc", x"cb",
    x"0f", x"19", x"1e", x"19", x"f9", x"01", x"19", x"ed",
    x"db", x"d3", x"21", x"11", x"1f", x"07", x"23", x"27",
    x"fe", x"21", x"d3", x"04", x"f8", x"f8", x"0a", x"f6",
    x"f6", x"03", x"f6", x"f4", x"ed", x"05", x"e2", x"11",
    x"2e", x"1f", x"03", x"18", x"20", x"fe", x"25", x"19",
    x"19", x"e3", x"e7", x"0c", x"1b", x"2a", x"b0", x"ed",
    x"d3", x"f9", x"15", x"20", x"16", x"f7", x"c1", x"c2",
    x"fa", x"28", x"03", x"06", x"2c", x"e1", x"04", x"7a",
    x"2c", x"24", x"f3", x"25", x"f5", x"27", x"fe", x"03",
    x"07", x"2b", x"12", x"36", x"1e", x"2e", x"23", x"06",
    x"ef", x"e6", x"17", x"ee", x"e9", x"3d", x"fd", x"df",
    x"8b", x"07", x"c3", x"43", x"50", x"e2", x"24", x"56",
    x"16", x"b9", x"27", x"05", x"04", x"f9", x"00", x"ff",
    x"04", x"01", x"00", x"01", x"02", x"1f", x"21", x"3a",
    x"ee", x"32", x"2e", x"e8", x"14", x"f4", x"69", x"ac",
    x"ba", x"f1", x"b1", x"26", x"df", x"f1", x"12", x"56",
    x"d8", x"dc", x"01", x"e7", x"04", x"ec", x"2d", x"16",
    x"00", x"ff", x"04", x"04", x"02", x"fc", x"fd", x"fc",
    x"01", x"ce", x"81", x"65", x"cd", x"0f", x"1d", x"0c",
    x"1c", x"09", x"21", x"00", x"ee", x"45", x"1c", x"37",
    x"ec", x"cd", x"e8", x"b1", x"d9", x"e7", x"43", x"10",
    x"f9", x"02", x"f1", x"96", x"b7", x"ef", x"c9", x"c0",
    x"21", x"37", x"09", x"1c", x"d2", x"09", x"ff", x"bb",
    x"1b", x"08", x"14", x"dc", x"e3", x"ed", x"cd", x"32",
    x"e9", x"14", x"0e", x"e5", x"ea", x"fa", x"03", x"dc",
    x"fa", x"02", x"1b", x"14", x"fe", x"df", x"f4", x"fe",
    x"03", x"03", x"01", x"07", x"03", x"fb", x"fe", x"00",
    x"fd", x"02", x"08", x"ff", x"00", x"06", x"06", x"01",
    x"08", x"fd", x"11", x"0f", x"19", x"ed", x"ec", x"be",
    x"9e", x"b5", x"ea", x"56", x"41", x"27", x"39", x"0f",
    x"5b", x"5b", x"2b", x"40", x"f3", x"ed", x"15", x"fc",
    x"15", x"0d", x"11", x"44", x"18", x"09", x"f6", x"0c",
    x"eb", x"16", x"fa", x"03", x"12", x"b1", x"a1", x"13",
    x"14", x"0d", x"fb", x"13", x"32", x"2a", x"26", x"0f",
    x"f6", x"cb", x"08", x"ed", x"01", x"4b", x"17", x"15",
    x"2f", x"1d", x"c8", x"36", x"c3", x"e8", x"f6", x"db",
    x"0d", x"2d", x"f8", x"04", x"de", x"d5", x"11", x"b7",
    x"ed", x"bd", x"0d", x"f1", x"98", x"e1", x"04", x"1b",
    x"c6", x"2f", x"ed", x"31", x"0a", x"fe", x"18", x"ef",
    x"e1", x"fa", x"9f", x"74", x"20", x"16", x"fe", x"4e",
    x"f0", x"f1", x"f7", x"ea", x"02", x"21", x"26", x"14",
    x"65", x"10", x"f7", x"02", x"fa", x"ea", x"37", x"f9",
    x"cd", x"18", x"ef", x"db", x"0f", x"de", x"d0", x"2a",
    x"04", x"09", x"2d", x"05", x"f0", x"17", x"c4", x"dd",
    x"2a", x"07", x"d7", x"31", x"4a", x"32", x"fe", x"50",
    x"56", x"08", x"2f", x"32", x"c1", x"fd", x"01", x"5a",
    x"1e", x"14", x"03", x"02", x"fc", x"f3", x"d9", x"e5",
    x"08", x"f4", x"d1", x"e3", x"cd", x"fe", x"db", x"ad",
    x"eb", x"0d", x"fc", x"fe", x"2a", x"e0", x"ee", x"09",
    x"1a", x"08", x"3c", x"21", x"44", x"f9", x"20", x"f3",
    x"bd", x"e1", x"08", x"db", x"ba", x"9e", x"2c", x"0a",
    x"24", x"cf", x"ff", x"10", x"ce", x"14", x"fb", x"26",
    x"0e", x"cd", x"07", x"18", x"22", x"f1", x"e9", x"07",
    x"23", x"37", x"0b", x"3b", x"42", x"51", x"06", x"40",
    x"48", x"ed", x"ce", x"e5", x"e5", x"ba", x"d7", x"57",
    x"3c", x"f7", x"35", x"fc", x"ec", x"d7", x"15", x"e9",
    x"51", x"3b", x"13", x"2c", x"0a", x"f1", x"16", x"ca",
    x"05", x"26", x"5d", x"59", x"38", x"f3", x"24", x"ed",
    x"13", x"fe", x"14", x"0f", x"0f", x"e9", x"d3", x"da",
    x"1f", x"e4", x"cd", x"09", x"23", x"49", x"ec", x"96",
    x"dd", x"16", x"b6", x"c8", x"18", x"e5", x"b8", x"09",
    x"87", x"86", x"15", x"d4", x"b8", x"17", x"d9", x"c8",
    x"0b", x"0a", x"f6", x"ef", x"09", x"ff", x"08", x"f5",
    x"0e", x"00", x"03", x"02", x"fd", x"ff", x"ff", x"03",
    x"01", x"fd", x"cf", x"a0", x"ed", x"c8", x"b5", x"e5",
    x"d1", x"b9", x"cb", x"19", x"0f", x"ef", x"e8", x"08",
    x"07", x"4f", x"0c", x"ed", x"f7", x"0c", x"ed", x"fa",
    x"df", x"fc", x"e9", x"03", x"10", x"bf", x"ef", x"ee",
    x"e3", x"fc", x"01", x"a4", x"b7", x"f1", x"f5", x"f0",
    x"ed", x"ec", x"f2", x"e3", x"e8", x"f7", x"0b", x"1e",
    x"2d", x"2a", x"2c", x"16", x"17", x"28", x"2b", x"40",
    x"4c", x"fd", x"16", x"03", x"0c", x"1d", x"3b", x"0b",
    x"33", x"e2", x"e0", x"e4", x"dc", x"d9", x"e1", x"c7",
    x"ef", x"1e", x"11", x"1b", x"e3", x"fb", x"16", x"16",
    x"b9", x"f5", x"2c", x"f8", x"04", x"ff", x"02", x"05",
    x"f9", x"00", x"ff", x"01", x"ed", x"df", x"cd", x"f8",
    x"eb", x"e9", x"ff", x"25", x"22", x"1c", x"2f", x"36",
    x"18", x"2b", x"13", x"cf", x"06", x"c1", x"e4", x"06",
    x"e8", x"1b", x"00", x"e4", x"07", x"0e", x"49", x"33",
    x"06", x"1b", x"0e", x"fe", x"00", x"ce", x"f1", x"19",
    x"0d", x"d8", x"ba", x"08", x"36", x"26", x"e1", x"f8",
    x"11", x"12", x"14", x"0f", x"02", x"ed", x"09", x"2c",
    x"4b", x"f6", x"f0", x"fd", x"e6", x"fc", x"cc", x"e9",
    x"d5", x"e2", x"fd", x"f1", x"08", x"24", x"35", x"00",
    x"02", x"0d", x"39", x"38", x"fc", x"fb", x"f8", x"f9",
    x"fa", x"f8", x"f9", x"fc", x"01", x"ec", x"fd", x"c5",
    x"bd", x"c2", x"d3", x"fe", x"ec", x"c5", x"0d", x"da",
    x"cd", x"42", x"fb", x"e5", x"1f", x"0b", x"fb", x"17",
    x"27", x"30", x"c0", x"ff", x"1b", x"e3", x"ef", x"0a",
    x"04", x"02", x"00", x"ff", x"00", x"ff", x"fb", x"02",
    x"03", x"0c", x"30", x"03", x"0f", x"37", x"31", x"01",
    x"09", x"16", x"3a", x"03", x"27", x"fe", x"10", x"16",
    x"d3", x"22", x"47", x"3b", x"23", x"16", x"6a", x"14",
    x"eb", x"4d", x"6d", x"62", x"d9", x"c5", x"27", x"e5",
    x"d2", x"e7", x"d6", x"d1", x"ea", x"46", x"47", x"44",
    x"0e", x"35", x"60", x"07", x"32", x"5e", x"00", x"d9",
    x"eb", x"03", x"e9", x"d8", x"e3", x"cd", x"d9", x"e0",
    x"cb", x"00", x"0e", x"cc", x"f1", x"17", x"e3", x"c6",
    x"ff", x"05", x"fb", x"01", x"fe", x"fb", x"00", x"01",
    x"fe", x"fa", x"01", x"f9", x"00", x"fc", x"fa", x"fc",
    x"fd", x"02", x"26", x"25", x"15", x"ff", x"fa", x"cf",
    x"11", x"ea", x"1b", x"e3", x"e1", x"d2", x"05", x"10",
    x"06", x"e0", x"ed", x"07", x"f8", x"eb", x"e1", x"df",
    x"d3", x"f5", x"b2", x"07", x"dc", x"07", x"f1", x"e7",
    x"10", x"0f", x"fe", x"cb", x"de", x"fd", x"dc", x"de",
    x"cc", x"a5", x"d5", x"b9", x"c9", x"bb", x"da", x"20",
    x"29", x"10", x"04", x"07", x"f6", x"a6", x"f1", x"e1",
    x"52", x"35", x"f7", x"16", x"f2", x"ee", x"fa", x"f6",
    x"0b", x"bb", x"0e", x"00", x"dc", x"0c", x"f5", x"03",
    x"0b", x"1f", x"c2", x"e6", x"0d", x"c1", x"b9", x"cb",
    x"ff", x"d4", x"96", x"ee", x"f0", x"ee", x"cd", x"e1",
    x"e9", x"dc", x"b2", x"b5", x"1e", x"38", x"2b", x"05",
    x"2e", x"33", x"19", x"2b", x"00", x"15", x"47", x"fb",
    x"fd", x"04", x"f3", x"e1", x"38", x"52", x"43", x"1c",
    x"ab", x"fe", x"49", x"3a", x"eb", x"d4", x"f4", x"49",
    x"2b", x"f9", x"e7", x"0e", x"07", x"fb", x"16", x"e8",
    x"0f", x"ff", x"f3", x"17", x"19", x"25", x"ff", x"0b",
    x"27", x"1d", x"d3", x"a5", x"24", x"ee", x"e5", x"1b",
    x"f4", x"d5", x"13", x"f4", x"e3", x"d0", x"ea", x"de",
    x"d9", x"cd", x"dd", x"24", x"0f", x"0a", x"e6", x"b5",
    x"f0", x"d9", x"ee", x"ea", x"32", x"d7", x"f9", x"00",
    x"ea", x"0e", x"f1", x"fb", x"d9", x"f6", x"21", x"04",
    x"00", x"08", x"1a", x"fd", x"00", x"f3", x"8d", x"cb",
    x"f5", x"92", x"c4", x"cc", x"56", x"31", x"3f", x"f3",
    x"e5", x"e1", x"49", x"2c", x"07", x"1b", x"fe", x"e9",
    x"19", x"d2", x"c5", x"30", x"06", x"ef", x"f6", x"dd",
    x"bd", x"0c", x"46", x"52", x"09", x"08", x"3d", x"c2",
    x"f2", x"fe", x"0c", x"0b", x"ea", x"3d", x"08", x"11",
    x"26", x"3a", x"18", x"dd", x"c9", x"e7", x"c8", x"df",
    x"14", x"fe", x"1c", x"2f", x"39", x"1a", x"cd", x"01",
    x"f6", x"f1", x"10", x"f4", x"04", x"a0", x"7b", x"11",
    x"ad", x"ae", x"c8", x"03", x"18", x"26", x"a5", x"1b",
    x"1f", x"5b", x"34", x"1c", x"36", x"29", x"33", x"17",
    x"08", x"1e", x"e7", x"01", x"30", x"31", x"0a", x"1d",
    x"f0", x"cc", x"f6", x"48", x"19", x"24", x"34", x"f4",
    x"08", x"fd", x"fe", x"03", x"04", x"fc", x"02", x"ff",
    x"05", x"fc", x"fa", x"fd", x"e0", x"6b", x"34", x"fa",
    x"05", x"03", x"13", x"04", x"dd", x"de", x"e0", x"dc",
    x"db", x"d9", x"03", x"dd", x"5b", x"a8", x"69", x"a1",
    x"da", x"1b", x"f6", x"14", x"13", x"3b", x"27", x"4d",
    x"19", x"ff", x"18", x"fe", x"f4", x"ea", x"eb", x"da",
    x"b9", x"01", x"1b", x"12", x"13", x"04", x"de", x"c0",
    x"a1", x"e4", x"f7", x"fd", x"26", x"48", x"08", x"fe",
    x"e0", x"7c", x"55", x"dc", x"c2", x"ca", x"70", x"2e",
    x"31", x"3e", x"33", x"18", x"e3", x"16", x"3a", x"01",
    x"2b", x"26", x"07", x"24", x"2f", x"2f", x"fe", x"0b",
    x"b0", x"70", x"b7", x"02", x"fc", x"04", x"03", x"0a",
    x"05", x"f9", x"ff", x"08", x"29", x"eb", x"63", x"1e",
    x"00", x"22", x"fc", x"f2", x"fe", x"e8", x"cb", x"c3",
    x"03", x"0d", x"fd", x"cc", x"0a", x"52", x"ec", x"cc",
    x"79", x"1d", x"21", x"19", x"39", x"12", x"1d", x"08",
    x"29", x"10", x"20", x"1e", x"0f", x"2e", x"1b", x"fd",
    x"e5", x"e3", x"a9", x"06", x"e6", x"15", x"e7", x"16",
    x"5a", x"13", x"fa", x"17", x"ad", x"f2", x"15", x"0a",
    x"03", x"1c", x"2f", x"19", x"0b", x"0f", x"14", x"26",
    x"03", x"1b", x"1c", x"53", x"c1", x"11", x"e6", x"f3",
    x"ea", x"08", x"e7", x"dd", x"03", x"0c", x"0a", x"04",
    x"0d", x"0a", x"07", x"0f", x"0a", x"c2", x"e7", x"dd",
    x"f6", x"db", x"09", x"5e", x"15", x"10", x"ce", x"e7",
    x"d5", x"17", x"1f", x"11", x"61", x"30", x"14", x"76",
    x"9c", x"df", x"e6", x"13", x"24", x"15", x"6c", x"50",
    x"01", x"05", x"05", x"fd", x"02", x"fb", x"03", x"02",
    x"fc", x"16", x"21", x"01", x"f3", x"f8", x"f2", x"32",
    x"09", x"08", x"50", x"55", x"19", x"02", x"f9", x"0b",
    x"1f", x"0a", x"f2", x"ed", x"00", x"cd", x"09", x"dd",
    x"cb", x"39", x"d1", x"dd", x"0a", x"18", x"b7", x"cc",
    x"02", x"de", x"ed", x"de", x"ef", x"7f", x"4e", x"b9",
    x"e3", x"fe", x"e6", x"17", x"0d", x"fa", x"4f", x"1e",
    x"b8", x"b7", x"cc", x"fb", x"ee", x"e3", x"ef", x"f8",
    x"fd", x"0a", x"d2", x"07", x"01", x"fa", x"08", x"12",
    x"fa", x"02", x"04", x"fd", x"fe", x"00", x"01", x"03",
    x"ff", x"04", x"08", x"03", x"05", x"03", x"05", x"00",
    x"04", x"01", x"bf", x"a2", x"4b", x"0c", x"10", x"12",
    x"d2", x"e8", x"f8", x"a7", x"af", x"dd", x"ea", x"dd",
    x"3e", x"f6", x"32", x"53", x"23", x"44", x"27", x"b9",
    x"12", x"14", x"da", x"e3", x"14", x"0b", x"ed", x"34",
    x"1b", x"12", x"0c", x"01", x"db", x"bf", x"3f", x"2d",
    x"36", x"36", x"35", x"0c", x"b2", x"f9", x"e6", x"ab",
    x"9b", x"94", x"cb", x"db", x"da", x"2e", x"14", x"29",
    x"0b", x"05", x"89", x"02", x"c7", x"df", x"24", x"0e",
    x"46", x"bf", x"eb", x"22", x"15", x"fd", x"f1", x"06",
    x"d0", x"ed", x"b3", x"28", x"e0", x"09", x"1d", x"11",
    x"41", x"2c", x"3a", x"15", x"2c", x"25", x"19", x"0f",
    x"17", x"02", x"00", x"d5", x"41", x"1e", x"1e", x"26",
    x"e0", x"01", x"e4", x"dc", x"f1", x"c3", x"45", x"39",
    x"e2", x"3b", x"18", x"22", x"05", x"f0", x"22", x"e7",
    x"d6", x"60", x"0f", x"f3", x"19", x"f9", x"ef", x"fd",
    x"12", x"1c", x"ca", x"ef", x"16", x"1b", x"04", x"f3",
    x"02", x"fd", x"fc", x"fe", x"01", x"fd", x"fc", x"fe",
    x"ff", x"fc", x"fa", x"fd", x"f8", x"fd", x"f9", x"02",
    x"fc", x"f7", x"fe", x"04", x"01", x"fa", x"f9", x"fc",
    x"02", x"01", x"fd", x"f8", x"f8", x"00", x"f8", x"fd",
    x"fd", x"04", x"fe", x"04", x"00", x"04", x"ff", x"f7",
    x"00", x"fc", x"00", x"fe", x"fb", x"01", x"01", x"03",
    x"ff", x"fd", x"ff", x"f8", x"fe", x"01", x"fe", x"fe",
    x"01", x"03", x"ff", x"fc", x"02", x"f9", x"fd", x"fc",
    x"fd", x"fd", x"ff", x"fb", x"fb", x"00", x"ff", x"fb",
    x"01", x"03", x"04", x"01", x"fd", x"03", x"fc", x"fa",
    x"00", x"ff", x"fe", x"f9", x"fb", x"fa", x"fd", x"fa",
    x"fa", x"f9", x"fb", x"fd", x"f9", x"fe", x"fe", x"f9",
    x"04", x"02", x"f7", x"01", x"01", x"fa", x"03", x"04",
    x"fd", x"02", x"fc", x"ff", x"01", x"01", x"f7", x"02",
    x"05", x"fc", x"fb", x"fc", x"00", x"fc", x"01", x"fd",
    x"fa", x"f7", x"01", x"f7", x"f9", x"04", x"fc", x"fd",
    x"fb", x"02", x"f9", x"01", x"fd", x"fd", x"fc", x"04",
    x"f7", x"04", x"f8", x"fa", x"04", x"00", x"f8", x"fe",
    x"02", x"fd", x"00", x"fd", x"fb", x"fa", x"fa", x"fd",
    x"fc", x"00", x"fd", x"fc", x"02", x"fd", x"03", x"00",
    x"02", x"02", x"fe", x"ff", x"ff", x"fb", x"ff", x"fe",
    x"fb", x"fe", x"ff", x"fd", x"01", x"ff", x"fb", x"02",
    x"02", x"ff", x"ff", x"f8", x"00", x"fd", x"00", x"ff",
    x"fa", x"fe", x"01", x"fe", x"fd", x"04", x"01", x"00",
    x"fb", x"ff", x"fc", x"fd", x"fe", x"03", x"fe", x"fb",
    x"01", x"04", x"f8", x"fe", x"fe", x"fa", x"fb", x"02",
    x"00", x"04", x"ff", x"fd", x"fb", x"fe", x"f9", x"fc",
    x"00", x"00", x"01", x"ff", x"02", x"01", x"00", x"00",
    x"fa", x"fe", x"fa", x"03", x"01", x"00", x"fe", x"fe",
    x"00", x"fd", x"03", x"fe", x"fd", x"f9", x"01", x"fa",
    x"fd", x"ff", x"00", x"03", x"00", x"02", x"05", x"02",
    x"fc", x"fc", x"fb", x"fc", x"fc", x"fe", x"fd", x"fa",
    x"fa", x"ff", x"f9", x"f9", x"00", x"fe", x"fe", x"00",
    x"00", x"fb", x"02", x"02", x"fb", x"fb", x"fb", x"fd",
    x"03", x"f8", x"fc", x"01", x"ff", x"01", x"02", x"ff",
    x"ff", x"fe", x"00", x"ff", x"ff", x"fb", x"fc", x"fd",
    x"fd", x"fb", x"f8", x"fc", x"fa", x"fb", x"f9", x"f9",
    x"03", x"fc", x"fb", x"00", x"00", x"ff", x"f9", x"01",
    x"fc", x"fc", x"fe", x"fb", x"fe", x"fb", x"fd", x"fc",
    x"01", x"00", x"ff", x"f8", x"fc", x"fa", x"ff", x"ff",
    x"fa", x"fe", x"fe", x"fe", x"00", x"fc", x"fc", x"fd",
    x"05", x"fb", x"02", x"fe", x"fc", x"fb", x"fe", x"04",
    x"02", x"fd", x"00", x"ff", x"f8", x"f8", x"fb", x"03",
    x"fc", x"00", x"03", x"fe", x"04", x"f9", x"ff", x"fa",
    x"fb", x"fb", x"fd", x"fb", x"f9", x"f7", x"ff", x"04",
    x"fc", x"fb", x"fb", x"04", x"04", x"fd", x"04", x"fc",
    x"02", x"02", x"fd", x"fe", x"05", x"f9", x"00", x"fb",
    x"f9", x"fb", x"fa", x"02", x"02", x"fd", x"f9", x"f9",
    x"fb", x"fb", x"f9", x"04", x"fc", x"fc", x"fe", x"fb",
    x"fa", x"03", x"ff", x"00", x"fd", x"01", x"fd", x"fe",
    x"03", x"04", x"fd", x"fa", x"ff", x"03", x"fc", x"fa",
    x"00", x"01", x"fa", x"fe", x"f8", x"fe", x"01", x"fe",
    x"02", x"f9", x"03", x"ff", x"ff", x"01", x"fd", x"00",
    x"ff", x"02", x"f8", x"fa", x"f7", x"fd", x"01", x"fa",
    x"ff", x"01", x"03", x"01", x"00", x"ff", x"02", x"02",
    x"04", x"00", x"02", x"02", x"fc", x"04", x"00", x"fb",
    x"fe", x"05", x"f7", x"03", x"fd", x"01", x"fe", x"f9",
    x"00", x"ff", x"fd", x"00", x"fc", x"04", x"fa", x"f9",
    x"03", x"f8", x"fc", x"fa", x"04", x"fd", x"00", x"00",
    x"fd", x"00", x"ff", x"ff", x"03", x"fb", x"fd", x"fc",
    x"f8", x"f7", x"fd", x"fa", x"04", x"ff", x"ff", x"03",
    x"fc", x"f8", x"fc", x"f8", x"fe", x"01", x"fd", x"02",
    x"03", x"04", x"ff", x"05", x"ff", x"fe", x"01", x"f8",
    x"fd", x"fe", x"fd", x"f8", x"02", x"04", x"05", x"fe",
    x"f9", x"fa", x"f8", x"fa", x"fc", x"fb", x"f8", x"f9",
    x"fa", x"fb", x"ff", x"01", x"ff", x"04", x"02", x"fa",
    x"ff", x"ff", x"fb", x"01", x"fe", x"fd", x"f8", x"01",
    x"00", x"fc", x"00", x"fa", x"fb", x"00", x"fc", x"04",
    x"fe", x"00", x"fb", x"00", x"f7", x"f8", x"f8", x"fe",
    x"fa", x"fd", x"fa", x"00", x"f8", x"fe", x"02", x"f8",
    x"fc", x"fb", x"fb", x"f9", x"fa", x"f7", x"fc", x"01",
    x"ff", x"03", x"fc", x"ff", x"fe", x"fa", x"fe", x"01",
    x"29", x"18", x"1a", x"2a", x"33", x"69", x"15", x"2c",
    x"7a", x"0d", x"08", x"f3", x"23", x"04", x"05", x"04",
    x"f2", x"e4", x"3e", x"2a", x"16", x"2c", x"38", x"2e",
    x"e2", x"ef", x"fd", x"b8", x"97", x"cb", x"de", x"e8",
    x"e5", x"36", x"03", x"e5", x"11", x"fc", x"d3", x"3a",
    x"0f", x"f5", x"fb", x"e9", x"e0", x"24", x"e9", x"e5",
    x"f0", x"07", x"4d", x"e5", x"26", x"16", x"20", x"21",
    x"23", x"f9", x"e3", x"e9", x"cd", x"ca", x"cd", x"dc",
    x"11", x"47", x"08", x"f7", x"19", x"17", x"0c", x"ef",
    x"f9", x"f9", x"eb", x"07", x"ff", x"fb", x"21", x"1b",
    x"45", x"05", x"e4", x"ea", x"65", x"88", x"c9", x"a2",
    x"cc", x"ec", x"79", x"de", x"07", x"7c", x"26", x"ee",
    x"44", x"a5", x"fb", x"2d", x"1d", x"f6", x"f6", x"bc",
    x"c3", x"d7", x"9c", x"e6", x"d8", x"ff", x"02", x"42",
    x"18", x"15", x"f9", x"03", x"12", x"09", x"31", x"2e",
    x"10", x"08", x"bf", x"ee", x"d6", x"b8", x"33", x"0d",
    x"2d", x"d3", x"02", x"20", x"f4", x"f4", x"0b", x"18",
    x"03", x"40", x"e6", x"f5", x"f0", x"af", x"cc", x"f4",
    x"e2", x"df", x"f1", x"09", x"fa", x"e7", x"0d", x"f7",
    x"f6", x"fc", x"fe", x"06", x"fc", x"fb", x"05", x"05",
    x"fc", x"04", x"1b", x"e9", x"e4", x"ec", x"f8", x"06",
    x"f6", x"fd", x"04", x"f8", x"09", x"f6", x"ed", x"0e",
    x"de", x"16", x"86", x"0a", x"37", x"31", x"5b", x"cb",
    x"a5", x"9e", x"ea", x"de", x"ce", x"eb", x"fa", x"1d",
    x"f5", x"f6", x"f6", x"ee", x"e2", x"a4", x"1a", x"12",
    x"ea", x"0f", x"28", x"32", x"29", x"f7", x"1e", x"06",
    x"02", x"e3", x"44", x"17", x"13", x"14", x"15", x"25",
    x"62", x"0f", x"00", x"2d", x"19", x"f2", x"f9", x"18",
    x"ea", x"49", x"2e", x"10", x"e1", x"01", x"0a", x"e0",
    x"ef", x"e5", x"03", x"f9", x"10", x"28", x"18", x"e3",
    x"65", x"0e", x"17", x"ff", x"03", x"09", x"02", x"06",
    x"04", x"01", x"05", x"04", x"1a", x"c7", x"00", x"02",
    x"e1", x"d5", x"19", x"20", x"f7", x"f9", x"e0", x"0a",
    x"47", x"39", x"64", x"24", x"22", x"ec", x"16", x"ec",
    x"f1", x"c4", x"b6", x"b3", x"85", x"a3", x"bd", x"dc",
    x"ec", x"fb", x"00", x"e4", x"e4", x"30", x"0f", x"ec",
    x"27", x"00", x"15", x"46", x"23", x"20", x"17", x"f3",
    x"ce", x"10", x"f1", x"01", x"b5", x"a4", x"97", x"e2",
    x"f5", x"35", x"36", x"2b", x"0e", x"34", x"1b", x"29",
    x"fb", x"34", x"40", x"2a", x"26", x"f5", x"2a", x"ea",
    x"d8", x"22", x"a8", x"c1", x"03", x"0e", x"05", x"f8",
    x"07", x"12", x"06", x"0f", x"08", x"07", x"f8", x"f2",
    x"f2", x"20", x"f7", x"d1", x"cf", x"d1", x"6a", x"14",
    x"0f", x"67", x"1e", x"23", x"2d", x"24", x"06", x"1f",
    x"3a", x"4b", x"38", x"26", x"15", x"1c", x"13", x"03",
    x"00", x"00", x"ff", x"03", x"03", x"03", x"01", x"07",
    x"fe", x"f3", x"ec", x"e0", x"15", x"09", x"0e", x"cc",
    x"8c", x"dc", x"f9", x"d9", x"d9", x"0e", x"e5", x"cb",
    x"3c", x"e5", x"cf", x"15", x"d9", x"d9", x"23", x"d7",
    x"d3", x"e6", x"fe", x"0e", x"1c", x"25", x"33", x"33",
    x"4a", x"36", x"34", x"0f", x"0a", x"07", x"1d", x"0e",
    x"1d", x"02", x"f9", x"22", x"38", x"4f", x"05", x"25",
    x"06", x"ec", x"fb", x"2d", x"d4", x"0e", x"23", x"0d",
    x"4a", x"30", x"2b", x"49", x"7e", x"00", x"26", x"3e",
    x"06", x"01", x"fa", x"ff", x"fd", x"04", x"ff", x"05",
    x"01", x"fa", x"ff", x"08", x"04", x"f9", x"fa", x"02",
    x"fb", x"ff", x"3f", x"1b", x"2c", x"47", x"32", x"30",
    x"32", x"43", x"41", x"38", x"43", x"35", x"31", x"0f",
    x"00", x"fa", x"bf", x"c1", x"f3", x"09", x"19", x"fa",
    x"1f", x"22", x"d7", x"c1", x"ee", x"fe", x"f1", x"00",
    x"02", x"24", x"3d", x"12", x"21", x"62", x"70", x"50",
    x"1f", x"f8", x"ed", x"f0", x"2e", x"0a", x"0d", x"30",
    x"36", x"2a", x"0d", x"f7", x"fe", x"fc", x"f0", x"09",
    x"32", x"01", x"09", x"b9", x"cf", x"c1", x"19", x"b7",
    x"c6", x"ba", x"d2", x"fe", x"01", x"fe", x"de", x"1f",
    x"e6", x"f5", x"3a", x"20", x"1f", x"f7", x"0e", x"1a",
    x"cb", x"f3", x"0b", x"2e", x"0c", x"1a", x"2d", x"0f",
    x"22", x"14", x"31", x"09", x"2e", x"d6", x"e4", x"ee",
    x"e5", x"ec", x"d9", x"f3", x"03", x"b6", x"07", x"21",
    x"d8", x"ec", x"d8", x"cb", x"f0", x"c0", x"0f", x"f1",
    x"12", x"26", x"32", x"51", x"46", x"28", x"28", x"1d",
    x"4a", x"3a", x"e3", x"59", x"44", x"13", x"3a", x"86",
    x"2b", x"2f", x"70", x"3d", x"36", x"9a", x"01", x"e7",
    x"4c", x"e6", x"e6", x"90", x"14", x"05", x"f1", x"e0",
    x"16", x"27", x"af", x"a0", x"e3", x"b9", x"ed", x"c5",
    x"08", x"e1", x"f1", x"e4", x"04", x"0a", x"d6", x"bf",
    x"f6", x"e3", x"0f", x"e7", x"cf", x"de", x"ef", x"cb",
    x"c4", x"0a", x"de", x"cb", x"c9", x"e7", x"1a", x"07",
    x"fa", x"ff", x"3d", x"de", x"ff", x"fb", x"e9", x"22",
    x"e1", x"02", x"c4", x"e9", x"f0", x"05", x"0e", x"07",
    x"c7", x"e1", x"eb", x"05", x"31", x"ca", x"e1", x"f1",
    x"1f", x"36", x"03", x"0d", x"00", x"df", x"d0", x"eb",
    x"f8", x"ef", x"40", x"20", x"44", x"2c", x"35", x"10",
    x"19", x"35", x"d9", x"c1", x"b4", x"21", x"c7", x"db",
    x"f2", x"ff", x"ed", x"1d", x"e4", x"d5", x"1d", x"f7",
    x"ef", x"f0", x"d3", x"cc", x"06", x"e9", x"f4", x"22",
    x"20", x"43", x"09", x"c6", x"fb", x"e7", x"a3", x"1c",
    x"bf", x"8e", x"a9", x"01", x"ea", x"09", x"aa", x"fe",
    x"dc", x"f0", x"ff", x"df", x"20", x"1f", x"2f", x"02",
    x"e5", x"17", x"f6", x"13", x"f3", x"e6", x"ee", x"17",
    x"3e", x"26", x"10", x"d8", x"1b", x"13", x"e8", x"ef",
    x"27", x"fc", x"fb", x"02", x"fc", x"fe", x"fb", x"fd",
    x"03", x"fc", x"d6", x"aa", x"49", x"2c", x"e2", x"19",
    x"f7", x"ea", x"9e", x"fd", x"15", x"f6", x"f3", x"f1",
    x"f8", x"29", x"3f", x"26", x"f8", x"9d", x"c8", x"2a",
    x"1c", x"f7", x"01", x"0f", x"3d", x"05", x"fd", x"0b",
    x"16", x"fa", x"ed", x"2e", x"0c", x"fc", x"23", x"13",
    x"fc", x"04", x"1d", x"f1", x"e3", x"e8", x"28", x"0b",
    x"06", x"22", x"0a", x"00", x"c7", x"f9", x"b7", x"ea",
    x"d8", x"bf", x"df", x"3c", x"f8", x"f1", x"de", x"e8",
    x"fe", x"0e", x"c5", x"e1", x"2f", x"0c", x"17", x"1f",
    x"12", x"0b", x"07", x"15", x"1e", x"18", x"ea", x"05",
    x"bc", x"e6", x"f1", x"fb", x"02", x"03", x"05", x"00",
    x"04", x"fc", x"fb", x"fe", x"1f", x"03", x"15", x"f5",
    x"f2", x"d1", x"07", x"f4", x"d9", x"e6", x"c0", x"af",
    x"c1", x"a6", x"cf", x"08", x"16", x"18", x"e4", x"dd",
    x"9f", x"07", x"12", x"04", x"27", x"11", x"2c", x"fd",
    x"08", x"0d", x"0b", x"d5", x"e0", x"e8", x"ab", x"d1",
    x"13", x"95", x"ad", x"35", x"18", x"dc", x"fa", x"ef",
    x"f7", x"1d", x"0f", x"f2", x"41", x"0e", x"23", x"09",
    x"29", x"2b", x"f6", x"ea", x"d5", x"ed", x"f7", x"ec",
    x"cc", x"e4", x"b6", x"2c", x"84", x"24", x"73", x"43",
    x"ab", x"33", x"1f", x"10", x"02", x"ff", x"04", x"02",
    x"09", x"04", x"00", x"00", x"fc", x"f5", x"a7", x"67",
    x"1b", x"2d", x"d8", x"db", x"0c", x"20", x"00", x"d3",
    x"e2", x"51", x"e6", x"da", x"35", x"ed", x"0d", x"02",
    x"c5", x"aa", x"66", x"1a", x"2c", x"f2", x"f2", x"1f",
    x"02", x"01", x"fa", x"03", x"fe", x"03", x"fc", x"ff",
    x"01", x"18", x"da", x"06", x"f8", x"db", x"c3", x"33",
    x"1f", x"0e", x"ec", x"c5", x"08", x"23", x"02", x"c6",
    x"f7", x"0f", x"03", x"07", x"e0", x"fb", x"1d", x"04",
    x"d8", x"24", x"03", x"ef", x"df", x"b9", x"e0", x"00",
    x"eb", x"db", x"ce", x"ea", x"25", x"c3", x"80", x"ba",
    x"fe", x"15", x"e6", x"db", x"e4", x"15", x"9c", x"ef",
    x"56", x"16", x"df", x"18", x"1c", x"eb", x"93", x"13",
    x"50", x"1a", x"1e", x"31", x"0d", x"56", x"14", x"10",
    x"04", x"01", x"05", x"fd", x"01", x"01", x"03", x"03",
    x"01", x"fa", x"fd", x"fd", x"05", x"02", x"fb", x"03",
    x"05", x"03", x"51", x"27", x"24", x"14", x"1b", x"3e",
    x"d3", x"e0", x"0c", x"11", x"ec", x"5f", x"14", x"1d",
    x"af", x"01", x"38", x"5b", x"99", x"01", x"43", x"08",
    x"05", x"4d", x"12", x"32", x"1d", x"0b", x"21", x"09",
    x"f7", x"ed", x"ff", x"95", x"c4", x"e7", x"6e", x"48",
    x"04", x"4a", x"0f", x"51", x"26", x"f2", x"26", x"a8",
    x"e8", x"16", x"a4", x"f4", x"e5", x"f5", x"e3", x"23",
    x"ea", x"cf", x"a2", x"30", x"ee", x"d2", x"3f", x"cc",
    x"c5", x"21", x"00", x"e0", x"c7", x"f1", x"11", x"e0",
    x"09", x"1a", x"03", x"49", x"47", x"ff", x"ce", x"2e",
    x"13", x"1b", x"3d", x"34", x"e8", x"05", x"2a", x"20",
    x"33", x"e3", x"e1", x"b9", x"ef", x"e8", x"20", x"16",
    x"fd", x"1f", x"04", x"04", x"d4", x"0b", x"4e", x"20",
    x"20", x"ed", x"c6", x"e9", x"0c", x"09", x"04", x"03",
    x"fb", x"34", x"28", x"39", x"20", x"0c", x"d3", x"9b",
    x"b6", x"e5", x"d2", x"da", x"dc", x"e5", x"d2", x"e8",
    x"06", x"fc", x"0f", x"e5", x"ce", x"08", x"bf", x"d9",
    x"38", x"1a", x"f2", x"fe", x"e0", x"f3", x"06", x"fa",
    x"c3", x"02", x"ee", x"06", x"1e", x"ed", x"19", x"3f",
    x"dd", x"fc", x"0e", x"10", x"31", x"23", x"d9", x"bc",
    x"11", x"25", x"04", x"04", x"0c", x"1e", x"eb", x"ec",
    x"01", x"03", x"ae", x"b7", x"8b", x"e9", x"00", x"e5",
    x"ee", x"06", x"33", x"00", x"ff", x"51", x"ec", x"02",
    x"4c", x"f7", x"1b", x"32", x"c9", x"58", x"3a", x"03",
    x"09", x"f9", x"10", x"0e", x"34", x"3f", x"28", x"43",
    x"da", x"f1", x"01", x"0e", x"f0", x"30", x"0c", x"11",
    x"f3", x"24", x"16", x"e2", x"11", x"ed", x"c8", x"9f",
    x"b2", x"93", x"1c", x"0b", x"07", x"a4", x"ec", x"dc",
    x"e7", x"3a", x"f3", x"07", x"22", x"32", x"c0", x"00",
    x"17", x"c9", x"47", x"2f", x"0c", x"e8", x"ba", x"cc",
    x"b2", x"cc", x"aa", x"e0", x"03", x"f3", x"2a", x"1f",
    x"e1", x"f9", x"1b", x"f8", x"15", x"10", x"e4", x"af",
    x"bb", x"dc", x"fe", x"f9", x"0e", x"26", x"13", x"05",
    x"f3", x"0d", x"f3", x"d6", x"15", x"e6", x"b1", x"d0",
    x"05", x"05", x"d6", x"f2", x"eb", x"df", x"0c", x"0a",
    x"fa", x"05", x"02", x"03", x"00", x"fc", x"fc", x"04",
    x"01", x"02", x"ee", x"e8", x"b3", x"09", x"2f", x"07",
    x"31", x"3c", x"48", x"f8", x"1f", x"0b", x"17", x"17",
    x"e9", x"fc", x"b8", x"9f", x"18", x"23", x"21", x"0a",
    x"e4", x"db", x"06", x"cd", x"d5", x"22", x"12", x"dc",
    x"58", x"46", x"2b", x"36", x"20", x"f3", x"03", x"07",
    x"fa", x"f6", x"f5", x"ef", x"de", x"2f", x"2d", x"1f",
    x"1b", x"3a", x"10", x"09", x"25", x"c7", x"cf", x"e1",
    x"4b", x"1e", x"1e", x"18", x"d7", x"08", x"23", x"ee",
    x"ff", x"c7", x"ff", x"e9", x"cf", x"ba", x"ad", x"c7",
    x"c4", x"b4", x"02", x"05", x"00", x"16", x"1e", x"14",
    x"dc", x"f9", x"f9", x"fc", x"f9", x"fa", x"f6", x"fb",
    x"f7", x"f8", x"fa", x"f4", x"f1", x"b7", x"dc", x"08",
    x"13", x"16", x"12", x"e7", x"e3", x"13", x"03", x"07",
    x"df", x"ec", x"b6", x"e6", x"90", x"8f", x"e9", x"07",
    x"f6", x"f1", x"d8", x"c7", x"3a", x"01", x"da", x"04",
    x"05", x"e8", x"f3", x"f9", x"06", x"f4", x"14", x"21",
    x"f3", x"fd", x"f3", x"ef", x"f2", x"29", x"e3", x"3a",
    x"46", x"2e", x"1f", x"f3", x"0e", x"14", x"14", x"f8",
    x"ed", x"c2", x"1a", x"1d", x"e3", x"ea", x"d9", x"12",
    x"11", x"32", x"26", x"18", x"16", x"e9", x"18", x"f7",
    x"ed", x"be", x"d2", x"b2", x"fc", x"04", x"00", x"fe",
    x"f7", x"f5", x"f8", x"0a", x"fe", x"45", x"03", x"02",
    x"21", x"03", x"19", x"ff", x"e1", x"ef", x"f7", x"18",
    x"bf", x"b9", x"f6", x"f3", x"c3", x"3a", x"2a", x"f8",
    x"fd", x"21", x"00", x"20", x"09", x"c4", x"45", x"3a",
    x"fc", x"ff", x"fd", x"01", x"01", x"fc", x"fc", x"fb",
    x"04", x"ed", x"de", x"f2", x"0b", x"f4", x"06", x"1b",
    x"fa", x"e3", x"17", x"24", x"e3", x"4b", x"28", x"19",
    x"47", x"60", x"37", x"08", x"14", x"0a", x"30", x"e8",
    x"e7", x"03", x"ca", x"ad", x"1d", x"fd", x"1f", x"16",
    x"1e", x"10", x"f6", x"17", x"0b", x"db", x"0c", x"f2",
    x"1b", x"19", x"20", x"0b", x"ff", x"2c", x"e6", x"da",
    x"c4", x"d6", x"ed", x"e1", x"ee", x"e9", x"df", x"1c",
    x"29", x"d7", x"2c", x"25", x"e8", x"07", x"fb", x"18",
    x"02", x"ff", x"06", x"0a", x"ff", x"02", x"05", x"02",
    x"fd", x"ff", x"00", x"ff", x"ff", x"ff", x"04", x"fd",
    x"02", x"04", x"ea", x"cf", x"b2", x"c9", x"e0", x"f3",
    x"e4", x"bc", x"e5", x"0f", x"30", x"2d", x"fb", x"1a",
    x"1e", x"34", x"47", x"31", x"18", x"0c", x"fc", x"fb",
    x"1c", x"1a", x"22", x"09", x"20", x"f4", x"d8", x"e3",
    x"1d", x"23", x"25", x"29", x"d5", x"bb", x"e9", x"0b",
    x"04", x"12", x"24", x"14", x"31", x"38", x"4b", x"20",
    x"32", x"1f", x"32", x"00", x"1d", x"c7", x"15", x"2e",
    x"01", x"0f", x"f7", x"29", x"e7", x"fd", x"98", x"2e",
    x"05", x"f1", x"01", x"0a", x"f9", x"fd", x"c6", x"ad",
    x"bf", x"dc", x"db", x"f6", x"16", x"f5", x"cc", x"dd",
    x"11", x"f4", x"e6", x"ef", x"f1", x"f2", x"06", x"33",
    x"33", x"19", x"1e", x"35", x"3a", x"f4", x"c4", x"2f",
    x"16", x"ed", x"aa", x"9e", x"a3", x"07", x"fe", x"03",
    x"1d", x"ec", x"cd", x"d8", x"77", x"81", x"ea", x"ce",
    x"d4", x"05", x"0f", x"0b", x"25", x"d7", x"f1", x"12",
    x"11", x"0a", x"14", x"ee", x"e9", x"de", x"12", x"f0",
    x"2a", x"17", x"fa", x"21", x"19", x"28", x"09", x"0c",
    x"39", x"d7", x"a9", x"11", x"f8", x"d4", x"20", x"c2",
    x"f1", x"28", x"f0", x"e5", x"e5", x"02", x"ea", x"07",
    x"18", x"12", x"32", x"ee", x"b9", x"c4", x"04", x"f7",
    x"c3", x"ea", x"0d", x"c6", x"b3", x"87", x"ba", x"dc",
    x"eb", x"1b", x"fe", x"12", x"25", x"1d", x"e5", x"49",
    x"0f", x"9a", x"e7", x"f7", x"b8", x"f9", x"02", x"fe",
    x"25", x"2e", x"ea", x"fa", x"fc", x"17", x"02", x"00",
    x"06", x"12", x"15", x"e8", x"04", x"2f", x"0e", x"f1",
    x"d7", x"dd", x"ff", x"e0", x"dd", x"17", x"ea", x"d9",
    x"16", x"05", x"c8", x"05", x"10", x"ec", x"e0", x"f0",
    x"eb", x"fc", x"39", x"ce", x"df", x"14", x"ec", x"08",
    x"21", x"51", x"3d", x"34", x"51", x"18", x"54", x"4f",
    x"06", x"33", x"00", x"f2", x"00", x"06", x"3c", x"4e",
    x"02", x"18", x"3b", x"1d", x"22", x"cc", x"e2", x"a4",
    x"ee", x"fa", x"c2", x"18", x"35", x"04", x"fa", x"51",
    x"f0", x"23", x"16", x"0b", x"21", x"20", x"02", x"ee",
    x"06", x"33", x"1d", x"24", x"ec", x"30", x"24", x"eb",
    x"ba", x"f2", x"3d", x"1c", x"de", x"2f", x"27", x"fc",
    x"07", x"02", x"fd", x"02", x"02", x"05", x"04", x"fe",
    x"04", x"fc", x"ca", x"16", x"ee", x"fe", x"02", x"e8",
    x"e7", x"05", x"0b", x"ba", x"c7", x"f8", x"b0", x"b6",
    x"24", x"bc", x"ce", x"01", x"ee", x"f8", x"c3", x"d9",
    x"1b", x"c8", x"fb", x"fd", x"02", x"bd", x"bf", x"fa",
    x"bf", x"c1", x"25", x"c3", x"c5", x"2b", x"f0", x"10",
    x"1a", x"de", x"d5", x"1c", x"09", x"03", x"5b", x"c5",
    x"f8", x"03", x"11", x"fb", x"fa", x"fd", x"41", x"5d",
    x"50", x"4f", x"1a", x"58", x"04", x"1e", x"26", x"d6",
    x"0e", x"1c", x"06", x"ad", x"55", x"44", x"08", x"fd",
    x"31", x"16", x"c9", x"bb", x"d7", x"e4", x"f6", x"06",
    x"ba", x"00", x"03", x"fc", x"0c", x"03", x"f6", x"0d",
    x"01", x"f8", x"04", x"02", x"f4", x"f0", x"3a", x"f8",
    x"e6", x"fd", x"fd", x"e3", x"22", x"ff", x"e9", x"2a",
    x"21", x"18", x"45", x"cf", x"bb", x"02", x"f3", x"cc",
    x"ef", x"12", x"0e", x"08", x"34", x"fe", x"e7", x"c1",
    x"e7", x"05", x"fb", x"fc", x"e4", x"2a", x"fd", x"f0",
    x"50", x"69", x"74", x"36", x"59", x"44", x"1c", x"07",
    x"15", x"e4", x"cc", x"dd", x"e8", x"fc", x"db", x"f3",
    x"30", x"2e", x"2e", x"59", x"4b", x"5a", x"36", x"1c",
    x"34", x"48", x"52", x"22", x"03", x"11", x"e5", x"de",
    x"c4", x"c1", x"df", x"e7", x"f8", x"03", x"02", x"f1",
    x"04", x"0d", x"fb", x"04", x"06", x"f5", x"93", x"55",
    x"ec", x"c0", x"98", x"28", x"f3", x"b7", x"40", x"e8",
    x"1f", x"4f", x"16", x"1d", x"51", x"13", x"f4", x"3b",
    x"f8", x"03", x"00", x"e4", x"e6", x"26", x"02", x"e2",
    x"fe", x"fb", x"fe", x"fb", x"00", x"03", x"fe", x"04",
    x"05", x"ea", x"af", x"c7", x"b3", x"b8", x"d9", x"e4",
    x"be", x"de", x"f0", x"b1", x"be", x"e9", x"c1", x"f3",
    x"d4", x"a8", x"1e", x"1d", x"e5", x"d9", x"fd", x"ef",
    x"f3", x"32", x"06", x"15", x"af", x"bf", x"cf", x"ef",
    x"ce", x"aa", x"f2", x"ea", x"f7", x"df", x"fc", x"ff",
    x"f1", x"e7", x"e1", x"19", x"0d", x"fd", x"7c", x"d4",
    x"52", x"f7", x"c8", x"5d", x"13", x"19", x"15", x"82",
    x"a6", x"12", x"e2", x"eb", x"f6", x"fe", x"fb", x"07",
    x"06", x"fc", x"fa", x"f5", x"fd", x"04", x"03", x"ff",
    x"03", x"fc", x"00", x"04", x"06", x"ff", x"03", x"fe",
    x"02", x"00", x"ed", x"1f", x"27", x"8b", x"13", x"1a",
    x"1f", x"18", x"22", x"ee", x"34", x"0a", x"d6", x"fb",
    x"e7", x"f4", x"00", x"10", x"ce", x"cb", x"c1", x"f2",
    x"ea", x"be", x"ef", x"1c", x"c6", x"de", x"fd", x"25",
    x"dd", x"ec", x"24", x"a2", x"ff", x"4a", x"fe", x"20",
    x"2c", x"0c", x"13", x"10", x"ba", x"dd", x"0d", x"53",
    x"13", x"2e", x"73", x"34", x"19", x"16", x"25", x"22",
    x"27", x"2e", x"20", x"37", x"18", x"18", x"f7", x"02",
    x"cd", x"26", x"08", x"1a", x"df", x"e2", x"25", x"a7",
    x"f8", x"29", x"09", x"30", x"24", x"b3", x"11", x"11",
    x"96", x"f3", x"03", x"6e", x"0a", x"2b", x"f5", x"23",
    x"30", x"19", x"14", x"27", x"18", x"25", x"5f", x"d9",
    x"ca", x"25", x"cc", x"f1", x"4f", x"4f", x"dd", x"0e",
    x"8e", x"be", x"cb", x"75", x"f5", x"02", x"22", x"0f",
    x"33", x"2f", x"01", x"14", x"45", x"e8", x"16", x"a3",
    x"28", x"85", x"f1", x"09", x"2c", x"07", x"06", x"7f",
    x"0a", x"26", x"2c", x"f9", x"01", x"0b", x"0e", x"f6",
    x"0d", x"1e", x"00", x"b2", x"fd", x"00", x"f6", x"f7",
    x"26", x"45", x"ea", x"ec", x"fe", x"24", x"35", x"1f",
    x"03", x"64", x"28", x"ef", x"df", x"fa", x"0d", x"f8",
    x"27", x"eb", x"ff", x"28", x"0b", x"1a", x"f3", x"1b",
    x"f0", x"cb", x"ee", x"c3", x"c3", x"9d", x"d8", x"e8",
    x"ef", x"dc", x"13", x"ec", x"14", x"fb", x"68", x"fe",
    x"16", x"0c", x"eb", x"d8", x"dc", x"bb", x"d8", x"91",
    x"ca", x"e9", x"e3", x"aa", x"05", x"d4", x"e7", x"f6",
    x"fe", x"ea", x"f4", x"03", x"e8", x"e5", x"16", x"01",
    x"c7", x"cc", x"d8", x"05", x"eb", x"17", x"3a", x"f9",
    x"06", x"d6", x"2d", x"14", x"fd", x"d3", x"2d", x"13",
    x"2d", x"6e", x"2f", x"f3", x"18", x"28", x"b8", x"41",
    x"4a", x"00", x"26", x"05", x"44", x"27", x"21", x"f0",
    x"b2", x"0d", x"c0", x"e6", x"ea", x"1e", x"42", x"24",
    x"14", x"23", x"98", x"0e", x"0b", x"bb", x"e6", x"c3",
    x"73", x"cf", x"df", x"c7", x"9d", x"92", x"d1", x"53",
    x"5d", x"19", x"27", x"41", x"25", x"17", x"45", x"e1",
    x"aa", x"e8", x"e7", x"fc", x"0b", x"2b", x"22", x"0e",
    x"39", x"fe", x"02", x"fc", x"ff", x"02", x"01", x"05",
    x"fe", x"03", x"d6", x"98", x"e0", x"c8", x"da", x"eb",
    x"16", x"0c", x"fa", x"d8", x"da", x"df", x"ff", x"05",
    x"c5", x"0e", x"b7", x"df", x"08", x"2e", x"16", x"eb",
    x"36", x"01", x"05", x"da", x"f9", x"f7", x"ea", x"09",
    x"28", x"17", x"0a", x"55", x"2d", x"a1", x"ce", x"16",
    x"21", x"11", x"2b", x"25", x"20", x"2b", x"61", x"f3",
    x"2f", x"15", x"ff", x"10", x"cc", x"0a", x"3d", x"10",
    x"10", x"37", x"13", x"e1", x"51", x"ff", x"05", x"00",
    x"fd", x"1b", x"3e", x"0b", x"ea", x"22", x"06", x"c4",
    x"0f", x"27", x"25", x"ff", x"c8", x"e4", x"c4", x"c7",
    x"06", x"d8", x"8f", x"00", x"fd", x"00", x"06", x"00",
    x"fc", x"00", x"00", x"05", x"c2", x"c3", x"d6", x"0d",
    x"cb", x"e0", x"fb", x"01", x"fa", x"1c", x"27", x"63",
    x"1c", x"3b", x"5b", x"24", x"39", x"12", x"f6", x"f0",
    x"c8", x"fd", x"fb", x"de", x"00", x"d7", x"e9", x"96",
    x"af", x"d9", x"ee", x"87", x"99", x"d9", x"b4", x"6d",
    x"2d", x"18", x"39", x"08", x"1b", x"28", x"da", x"e5",
    x"f6", x"84", x"fa", x"d7", x"e7", x"00", x"cf", x"0d",
    x"e7", x"8b", x"15", x"d6", x"ed", x"d3", x"e3", x"f1",
    x"cd", x"ef", x"29", x"17", x"16", x"e4", x"e0", x"d3",
    x"ac", x"fd", x"bd", x"c4", x"06", x"0b", x"06", x"ff",
    x"fb", x"fb", x"06", x"03", x"05", x"12", x"0d", x"f5",
    x"4e", x"23", x"fa", x"05", x"e7", x"0b", x"f2", x"55",
    x"21", x"49", x"30", x"18", x"3e", x"fd", x"09", x"85",
    x"ff", x"f8", x"06", x"2b", x"32", x"ff", x"fe", x"00",
    x"fc", x"01", x"fe", x"04", x"04", x"04", x"03", x"02",
    x"fb", x"06", x"f7", x"cf", x"ef", x"f1", x"ff", x"04",
    x"f2", x"e9", x"14", x"56", x"e2", x"42", x"18", x"f5",
    x"27", x"c8", x"ba", x"33", x"eb", x"d7", x"bd", x"dc",
    x"ba", x"0f", x"e2", x"d3", x"15", x"4a", x"35", x"4a",
    x"3f", x"02", x"f0", x"14", x"15", x"c4", x"1b", x"09",
    x"11", x"f3", x"d8", x"cd", x"e3", x"d1", x"b6", x"d5",
    x"d9", x"d0", x"1a", x"10", x"0a", x"2d", x"07", x"d1",
    x"c5", x"d5", x"e4", x"e8", x"e4", x"04", x"21", x"ff",
    x"fc", x"fc", x"01", x"04", x"fc", x"01", x"00", x"05",
    x"04", x"fb", x"00", x"03", x"00", x"04", x"04", x"05",
    x"fd", x"ff", x"c0", x"00", x"e2", x"f8", x"0c", x"fd",
    x"e6", x"fe", x"47", x"fa", x"0f", x"f8", x"f7", x"f7",
    x"b9", x"da", x"db", x"c9", x"b7", x"bd", x"dd", x"de",
    x"dd", x"0c", x"09", x"0e", x"e9", x"1a", x"b5", x"f4",
    x"fb", x"c3", x"de", x"08", x"e4", x"f5", x"80", x"06",
    x"03", x"bb", x"15", x"1b", x"f9", x"10", x"00", x"da",
    x"fe", x"0a", x"3a", x"1d", x"f1", x"3f", x"fb", x"ed",
    x"f1", x"0b", x"14", x"ea", x"2c", x"14", x"13", x"2f",
    x"0e", x"ef", x"b2", x"a8", x"fd", x"dd", x"e0", x"e6",
    x"dc", x"f4", x"04", x"1b", x"30", x"1f", x"fb", x"21",
    x"d4", x"0d", x"03", x"a0", x"87", x"78", x"ea", x"fb",
    x"ca", x"0f", x"37", x"fe", x"17", x"ea", x"b8", x"04",
    x"27", x"fb", x"e5", x"ed", x"d6", x"c5", x"f1", x"f3",
    x"d5", x"e3", x"b5", x"fa", x"e2", x"f5", x"c3", x"b8",
    x"be", x"90", x"ff", x"12", x"bd", x"16", x"19", x"d5",
    x"03", x"03", x"e3", x"f6", x"17", x"ee", x"0b", x"13",
    x"37", x"c8", x"58", x"29", x"21", x"26", x"20", x"56",
    x"d2", x"02", x"0e", x"46", x"e1", x"05", x"16", x"fd",
    x"f2", x"d9", x"c8", x"c0", x"a7", x"c6", x"bc", x"b5",
    x"00", x"ef", x"ef", x"fb", x"01", x"15", x"ba", x"d8",
    x"10", x"ea", x"d0", x"03", x"ef", x"1d", x"18", x"e8",
    x"f7", x"04", x"fd", x"05", x"f0", x"e8", x"fa", x"1f",
    x"c2", x"ff", x"1a", x"ec", x"d8", x"ec", x"15", x"eb",
    x"db", x"03", x"e9", x"bc", x"23", x"22", x"dc", x"83",
    x"43", x"93", x"2e", x"1d", x"36", x"0c", x"17", x"09",
    x"35", x"3a", x"dc", x"2f", x"25", x"25", x"16", x"18",
    x"3c", x"e7", x"1a", x"19", x"dc", x"dd", x"db", x"ce",
    x"08", x"ff", x"19", x"d4", x"e5", x"ee", x"ee", x"ff",
    x"10", x"38", x"31", x"c3", x"d0", x"e2", x"98", x"e9",
    x"e0", x"ee", x"01", x"16", x"65", x"17", x"f1", x"1a",
    x"14", x"21", x"26", x"09", x"e2", x"a8", x"17", x"81",
    x"ae", x"af", x"b4", x"f0", x"e7", x"d1", x"44", x"e3",
    x"02", x"2e", x"e8", x"cc", x"14", x"ec", x"b4", x"ee",
    x"ad", x"e4", x"08", x"cc", x"e5", x"f0", x"fe", x"d8",
    x"25", x"61", x"3e", x"3e", x"55", x"67", x"f5", x"2c",
    x"58", x"01", x"01", x"01", x"fa", x"05", x"fc", x"02",
    x"ff", x"03", x"10", x"ee", x"34", x"11", x"f9", x"e3",
    x"f3", x"0e", x"fb", x"01", x"05", x"f6", x"f6", x"e9",
    x"08", x"14", x"d6", x"df", x"e8", x"02", x"12", x"11",
    x"e7", x"2d", x"0e", x"ca", x"e4", x"04", x"dd", x"0e",
    x"02", x"d3", x"f4", x"ea", x"f0", x"ec", x"28", x"f3",
    x"ec", x"2f", x"27", x"36", x"3b", x"1e", x"71", x"08",
    x"20", x"24", x"08", x"20", x"14", x"08", x"2e", x"20",
    x"19", x"02", x"e9", x"14", x"15", x"fe", x"32", x"1f",
    x"29", x"a6", x"e1", x"31", x"fe", x"0b", x"38", x"e5",
    x"26", x"46", x"0c", x"1e", x"ed", x"11", x"13", x"0b",
    x"fa", x"ff", x"29", x"01", x"f9", x"fa", x"ff", x"05",
    x"f6", x"f9", x"06", x"f7", x"19", x"22", x"1b", x"2c",
    x"11", x"11", x"13", x"1a", x"fd", x"1a", x"29", x"fb",
    x"ee", x"1d", x"39", x"e6", x"22", x"1e", x"a8", x"c6",
    x"cb", x"00", x"08", x"0d", x"01", x"f1", x"0f", x"36",
    x"20", x"ff", x"2b", x"20", x"4b", x"0e", x"fa", x"10",
    x"24", x"f5", x"06", x"ee", x"26", x"44", x"27", x"4f",
    x"42", x"fc", x"03", x"26", x"17", x"fe", x"4f", x"c6",
    x"27", x"fd", x"1e", x"ee", x"ec", x"bf", x"8a", x"a2",
    x"fa", x"c9", x"b3", x"1d", x"e8", x"ee", x"03", x"18",
    x"1e", x"a7", x"13", x"0d", x"ff", x"fe", x"ff", x"fd",
    x"00", x"f5", x"05", x"f8", x"f9", x"f4", x"ef", x"dd",
    x"bb", x"f2", x"07", x"e5", x"fd", x"29", x"08", x"fd",
    x"ff", x"11", x"07", x"da", x"4d", x"24", x"fc", x"01",
    x"ff", x"41", x"bf", x"dc", x"df", x"d0", x"03", x"ef",
    x"06", x"ff", x"ff", x"ff", x"fd", x"02", x"01", x"03",
    x"00", x"97", x"e9", x"1c", x"f5", x"02", x"fd", x"28",
    x"fc", x"00", x"21", x"ed", x"f0", x"1a", x"0a", x"f5",
    x"fe", x"2f", x"3a", x"fc", x"ec", x"2d", x"16", x"2c",
    x"04", x"23", x"0e", x"f8", x"a7", x"f3", x"f7", x"c0",
    x"ee", x"d3", x"e9", x"e6", x"f7", x"50", x"61", x"be",
    x"2e", x"3c", x"2c", x"32", x"58", x"2c", x"38", x"33",
    x"2a", x"1b", x"02", x"f9", x"db", x"f4", x"06", x"c3",
    x"ec", x"15", x"dc", x"aa", x"e9", x"03", x"ce", x"f7",
    x"04", x"fa", x"05", x"f5", x"fd", x"02", x"fc", x"fa",
    x"fd", x"fe", x"f8", x"03", x"01", x"00", x"01", x"fd",
    x"fb", x"01", x"24", x"25", x"43", x"f2", x"0e", x"14",
    x"13", x"18", x"1b", x"0f", x"14", x"f7", x"dc", x"3d",
    x"3a", x"fc", x"f2", x"f9", x"d5", x"db", x"02", x"cb",
    x"cc", x"ea", x"f6", x"e6", x"e7", x"ed", x"08", x"01",
    x"f9", x"06", x"3f", x"d4", x"00", x"da", x"04", x"cf",
    x"dd", x"f6", x"de", x"cf", x"d6", x"bf", x"c4", x"36",
    x"fc", x"d2", x"e4", x"ef", x"fb", x"1f", x"ff", x"3b",
    x"18", x"bf", x"af", x"16", x"e4", x"d4", x"12", x"3c",
    x"2f", x"e2", x"f5", x"22", x"dd", x"0b", x"25", x"b3",
    x"0a", x"10", x"04", x"c2", x"fd", x"03", x"af", x"9d",
    x"37", x"c7", x"cd", x"17", x"19", x"f5", x"fa", x"df",
    x"e7", x"ca", x"9b", x"d0", x"25", x"24", x"3d", x"4b",
    x"ed", x"fb", x"07", x"0f", x"e0", x"42", x"53", x"03",
    x"26", x"29", x"f1", x"e1", x"ea", x"d8", x"1c", x"f9",
    x"f1", x"09", x"01", x"f8", x"01", x"0c", x"01", x"0a",
    x"1c", x"ff", x"ff", x"f4", x"da", x"1a", x"c4", x"a7",
    x"15", x"f9", x"e2", x"04", x"14", x"14", x"09", x"fd",
    x"12", x"e8", x"0e", x"20", x"c1", x"db", x"ff", x"db",
    x"05", x"c5", x"f4", x"0b", x"19", x"d5", x"03", x"0e",
    x"cc", x"df", x"ef", x"0c", x"00", x"12", x"14", x"4f",
    x"10", x"11", x"2e", x"fe", x"0a", x"2a", x"f0", x"e0",
    x"eb", x"f8", x"90", x"88", x"a7", x"ba", x"d8", x"b8",
    x"c4", x"bc", x"b5", x"e3", x"cb", x"c4", x"e5", x"22",
    x"29", x"fd", x"f8", x"05", x"26", x"0a", x"06", x"ac",
    x"df", x"56", x"30", x"1d", x"0c", x"31", x"2e", x"14",
    x"e4", x"bd", x"e2", x"d5", x"fc", x"1d", x"ee", x"20",
    x"4e", x"b2", x"a0", x"ae", x"c4", x"a2", x"9e", x"12",
    x"fb", x"9b", x"13", x"11", x"da", x"fd", x"1b", x"e6",
    x"1f", x"1d", x"23", x"11", x"19", x"fd", x"1d", x"0b",
    x"07", x"43", x"32", x"36", x"2a", x"ba", x"d3", x"f2",
    x"bb", x"e0", x"e5", x"ab", x"bb", x"89", x"75", x"6b",
    x"ee", x"cd", x"a5", x"0f", x"f6", x"cd", x"0a", x"cb",
    x"72", x"e7", x"04", x"9f", x"0c", x"0b", x"08", x"e8",
    x"f2", x"eb", x"ca", x"d5", x"f3", x"c9", x"cd", x"e0",
    x"d6", x"0a", x"1d", x"d1", x"e4", x"fb", x"b2", x"cd",
    x"00", x"05", x"04", x"00", x"fd", x"01", x"fb", x"fe",
    x"fe", x"fc", x"c9", x"dc", x"b7", x"22", x"78", x"c4",
    x"33", x"49", x"24", x"b5", x"cd", x"cd", x"f1", x"15",
    x"0b", x"ea", x"b8", x"c2", x"d7", x"ed", x"cb", x"ef",
    x"e3", x"e9", x"12", x"1b", x"f1", x"ed", x"f5", x"f4",
    x"f5", x"ef", x"e9", x"e3", x"19", x"10", x"03", x"03",
    x"14", x"e4", x"06", x"0c", x"d5", x"cb", x"f5", x"1f",
    x"e9", x"bf", x"02", x"1e", x"12", x"ef", x"e8", x"f7",
    x"02", x"0b", x"fb", x"1a", x"39", x"12", x"ed", x"df",
    x"f0", x"13", x"f7", x"d8", x"e3", x"ec", x"02", x"fb",
    x"a9", x"ec", x"04", x"0e", x"06", x"0c", x"0f", x"20",
    x"bb", x"ed", x"f9", x"02", x"fe", x"02", x"fd", x"03",
    x"04", x"ff", x"fe", x"fc", x"f8", x"c8", x"ca", x"f4",
    x"13", x"e2", x"08", x"29", x"1e", x"0a", x"3e", x"02",
    x"2e", x"3f", x"28", x"e6", x"19", x"20", x"cb", x"b5",
    x"09", x"ec", x"ef", x"f3", x"11", x"19", x"fa", x"02",
    x"c8", x"e3", x"07", x"fa", x"ed", x"0b", x"49", x"3d",
    x"cc", x"eb", x"01", x"e0", x"08", x"12", x"28", x"37",
    x"2b", x"cd", x"e8", x"f4", x"d6", x"ea", x"1f", x"db",
    x"b6", x"e4", x"23", x"21", x"2c", x"1d", x"17", x"14",
    x"2d", x"45", x"22", x"df", x"da", x"d3", x"f3", x"00",
    x"05", x"5b", x"06", x"f6", x"07", x"0a", x"fc", x"00",
    x"10", x"07", x"07", x"0a", x"0d", x"05", x"1a", x"1b",
    x"e6", x"10", x"13", x"14", x"01", x"f1", x"f4", x"f9",
    x"ee", x"01", x"22", x"18", x"31", x"26", x"1c", x"f6",
    x"0e", x"f7", x"29", x"0a", x"05", x"2d", x"31", x"25",
    x"ff", x"00", x"05", x"fe", x"fb", x"01", x"04", x"03",
    x"01", x"16", x"0e", x"f6", x"00", x"ff", x"0a", x"11",
    x"02", x"c5", x"16", x"12", x"ca", x"33", x"4a", x"14",
    x"04", x"40", x"47", x"3b", x"0d", x"24", x"cf", x"35",
    x"2a", x"ef", x"01", x"e6", x"db", x"fe", x"25", x"82",
    x"bb", x"e5", x"d0", x"d0", x"ca", x"f4", x"f6", x"10",
    x"16", x"f8", x"f1", x"f0", x"e6", x"02", x"c0", x"f2",
    x"fe", x"dc", x"ee", x"f4", x"ca", x"da", x"f8", x"e6",
    x"a8", x"ff", x"d6", x"b7", x"bf", x"df", x"d5", x"c3",
    x"fe", x"04", x"fc", x"03", x"fd", x"fc", x"fe", x"00",
    x"fe", x"ff", x"02", x"ff", x"fb", x"00", x"02", x"fe",
    x"05", x"05", x"33", x"dd", x"dd", x"ea", x"f2", x"da",
    x"de", x"d3", x"e7", x"09", x"ea", x"f2", x"ff", x"31",
    x"08", x"17", x"0b", x"1b", x"c2", x"ee", x"d5", x"ca",
    x"b4", x"d0", x"ec", x"e5", x"ee", x"f9", x"ee", x"ee",
    x"36", x"24", x"18", x"20", x"3a", x"20", x"03", x"fa",
    x"f1", x"f4", x"bc", x"fe", x"f4", x"ec", x"e4", x"53",
    x"2d", x"f9", x"55", x"0a", x"ff", x"6d", x"2c", x"10",
    x"42", x"34", x"0a", x"1d", x"14", x"f7", x"0a", x"fb",
    x"13", x"25", x"fb", x"f4", x"26", x"ff", x"e2", x"ff",
    x"e1", x"e9", x"20", x"f3", x"12", x"0c", x"ff", x"f2",
    x"dc", x"fd", x"ea", x"e1", x"da", x"a6", x"03", x"dc",
    x"da", x"f3", x"f3", x"f4", x"fe", x"af", x"ff", x"54",
    x"32", x"16", x"f9", x"f8", x"fb", x"e4", x"01", x"f1",
    x"f7", x"fb", x"fa", x"ef", x"06", x"18", x"ef", x"e6",
    x"18", x"cd", x"e7", x"13", x"db", x"d0", x"e1", x"3d",
    x"65", x"20", x"2b", x"20", x"08", x"28", x"1a", x"25",
    x"1e", x"f6", x"2d", x"19", x"fe", x"0a", x"0e", x"04",
    x"d3", x"30", x"0d", x"f2", x"1a", x"00", x"07", x"e9",
    x"13", x"16", x"f2", x"f4", x"11", x"13", x"17", x"3b",
    x"f9", x"0b", x"13", x"f5", x"fa", x"08", x"18", x"4c",
    x"37", x"f5", x"f8", x"f1", x"25", x"fb", x"04", x"1c",
    x"f7", x"0e", x"f2", x"dc", x"fc", x"14", x"0a", x"fb",
    x"06", x"0a", x"16", x"00", x"37", x"35", x"0d", x"ea",
    x"f1", x"e9", x"fe", x"e9", x"da", x"da", x"bf", x"3f",
    x"5f", x"25", x"50", x"55", x"6b", x"2d", x"20", x"78",
    x"f4", x"00", x"24", x"0d", x"04", x"23", x"1f", x"1b",
    x"d4", x"db", x"e1", x"c0", x"d6", x"ed", x"cb", x"cb",
    x"da", x"c4", x"e8", x"1e", x"46", x"53", x"36", x"53",
    x"15", x"57", x"36", x"18", x"42", x"38", x"2e", x"14",
    x"0b", x"d2", x"0e", x"14", x"f4", x"fe", x"c2", x"46",
    x"0b", x"11", x"34", x"1d", x"3c", x"fe", x"f5", x"e7",
    x"f6", x"de", x"d6", x"d9", x"f3", x"12", x"17", x"3b",
    x"06", x"00", x"19", x"f7", x"f9", x"ca", x"c0", x"f1",
    x"34", x"fe", x"06", x"ef", x"e2", x"ee", x"ee", x"d5",
    x"18", x"ec", x"c8", x"e2", x"ea", x"b7", x"fa", x"23",
    x"23", x"05", x"02", x"fc", x"05", x"03", x"00", x"fc",
    x"05", x"fe", x"a6", x"d8", x"e5", x"f5", x"1b", x"22",
    x"08", x"21", x"0b", x"eb", x"dc", x"cc", x"bb", x"99",
    x"73", x"c9", x"aa", x"7c", x"15", x"f7", x"23", x"0a",
    x"03", x"cc", x"f6", x"06", x"e6", x"08", x"05", x"06",
    x"03", x"1e", x"16", x"52", x"48", x"2e", x"fa", x"19",
    x"23", x"13", x"19", x"39", x"4c", x"36", x"49", x"ea",
    x"2f", x"44", x"fb", x"22", x"2b", x"04", x"2d", x"25",
    x"2c", x"2d", x"0b", x"29", x"13", x"10", x"a7", x"12",
    x"ed", x"e7", x"0b", x"2d", x"c5", x"16", x"02", x"b5",
    x"fd", x"0d", x"f3", x"db", x"db", x"d3", x"01", x"ea",
    x"25", x"42", x"36", x"fb", x"fe", x"02", x"fc", x"fe",
    x"fd", x"04", x"fa", x"f5", x"10", x"43", x"4b", x"3b",
    x"48", x"2b", x"f5", x"12", x"02", x"22", x"52", x"4f",
    x"0e", x"2a", x"09", x"2f", x"0c", x"db", x"d5", x"e6",
    x"ea", x"f9", x"fc", x"0e", x"fb", x"d3", x"b4", x"3e",
    x"4c", x"26", x"3b", x"22", x"0f", x"31", x"2e", x"37",
    x"17", x"27", x"33", x"e8", x"01", x"f6", x"e6", x"f3",
    x"f8", x"ea", x"e6", x"f0", x"b2", x"0e", x"c0", x"18",
    x"15", x"13", x"1d", x"17", x"1d", x"31", x"04", x"ed",
    x"38", x"21", x"06", x"e7", x"0a", x"ee", x"21", x"da",
    x"d7", x"44", x"b3", x"a0", x"04", x"01", x"00", x"fe",
    x"fe", x"fd", x"0a", x"06", x"05", x"fb", x"f2", x"0c",
    x"22", x"eb", x"07", x"4c", x"22", x"fe", x"25", x"34",
    x"36", x"0c", x"05", x"0e", x"15", x"ed", x"c8", x"c4",
    x"fe", x"28", x"d5", x"fa", x"f9", x"dd", x"f7", x"df",
    x"00", x"fe", x"01", x"04", x"fd", x"05", x"02", x"06",
    x"02", x"f3", x"ec", x"d5", x"e7", x"cf", x"c3", x"f0",
    x"ad", x"8b", x"15", x"47", x"34", x"3d", x"54", x"26",
    x"3e", x"10", x"f3", x"1c", x"16", x"24", x"36", x"e8",
    x"e5", x"db", x"c7", x"d1", x"40", x"22", x"4c", x"11",
    x"fa", x"f8", x"08", x"24", x"11", x"5d", x"2d", x"21",
    x"05", x"f7", x"f0", x"fc", x"ea", x"ce", x"be", x"e0",
    x"f4", x"dc", x"cd", x"e8", x"df", x"f2", x"f5", x"a9",
    x"8f", x"bf", x"c2", x"cd", x"f9", x"f8", x"0b", x"22",
    x"03", x"00", x"fb", x"01", x"02", x"fc", x"01", x"00",
    x"05", x"f9", x"fd", x"03", x"04", x"02", x"03", x"04",
    x"06", x"00", x"07", x"d6", x"ef", x"0f", x"e5", x"ea",
    x"00", x"b9", x"cb", x"bf", x"fb", x"ff", x"be", x"f9",
    x"f2", x"cd", x"f0", x"e4", x"bc", x"b0", x"c9", x"e2",
    x"fc", x"04", x"19", x"31", x"12", x"f7", x"14", x"f4",
    x"d4", x"ec", x"0c", x"3b", x"6d", x"4b", x"c4", x"0c",
    x"0e", x"05", x"fc", x"18", x"1d", x"0e", x"02", x"1c",
    x"ed", x"f7", x"47", x"00", x"e4", x"0f", x"18", x"1e",
    x"21", x"29", x"0f", x"3e", x"59", x"4a", x"6b", x"fe",
    x"ee", x"e7", x"15", x"fa", x"a4", x"f9", x"20", x"fd",
    x"fb", x"00", x"e6", x"dd", x"fe", x"e4", x"e1", x"0b",
    x"e7", x"16", x"24", x"fd", x"11", x"e6", x"0b", x"08",
    x"09", x"39", x"2a", x"6e", x"00", x"fa", x"f6", x"fe",
    x"c7", x"db", x"01", x"d4", x"dc", x"db", x"e5", x"be",
    x"08", x"08", x"10", x"23", x"31", x"15", x"c1", x"d7",
    x"ac", x"16", x"0a", x"d9", x"31", x"43", x"47", x"3b",
    x"13", x"14", x"14", x"f0", x"f6", x"31", x"13", x"46",
    x"1c", x"1b", x"b9", x"2b", x"25", x"e5", x"01", x"09",
    x"21", x"1c", x"11", x"00", x"ca", x"29", x"37", x"b2",
    x"e3", x"f4", x"f4", x"fd", x"be", x"0e", x"96", x"9b",
    x"fb", x"fb", x"df", x"e9", x"af", x"e1", x"0c", x"c6",
    x"9d", x"f9", x"04", x"fd", x"d3", x"f0", x"e5", x"d6",
    x"d0", x"df", x"f7", x"b5", x"c4", x"bb", x"e6", x"1e",
    x"ec", x"0f", x"2c", x"b9", x"ce", x"c2", x"26", x"f5",
    x"30", x"32", x"05", x"eb", x"dc", x"8d", x"c6", x"83",
    x"d7", x"4b", x"e3", x"ee", x"22", x"1b", x"29", x"23",
    x"21", x"d8", x"0a", x"f7", x"e7", x"3b", x"05", x"24",
    x"59", x"88", x"cc", x"08", x"ec", x"f3", x"05", x"e6",
    x"26", x"25", x"5c", x"15", x"b9", x"09", x"8e", x"96",
    x"04", x"b3", x"e0", x"4c", x"3b", x"28", x"1a", x"11",
    x"c8", x"6f", x"43", x"14", x"dd", x"29", x"1a", x"56",
    x"1d", x"f6", x"e5", x"ed", x"e7", x"ac", x"b1", x"fb",
    x"ce", x"17", x"e1", x"05", x"0a", x"e5", x"de", x"f2",
    x"93", x"ed", x"02", x"01", x"0d", x"18", x"05", x"df",
    x"c4", x"10", x"ec", x"a1", x"c3", x"bf", x"90", x"cb",
    x"29", x"05", x"00", x"e4", x"f1", x"1b", x"d6", x"d9",
    x"22", x"ff", x"01", x"ff", x"fe", x"fc", x"01", x"03",
    x"ff", x"fe", x"c8", x"8b", x"b6", x"86", x"e3", x"f1",
    x"da", x"0a", x"22", x"53", x"3e", x"0b", x"e4", x"03",
    x"3d", x"30", x"31", x"28", x"29", x"3a", x"07", x"ea",
    x"c7", x"b2", x"de", x"dd", x"ef", x"eb", x"fa", x"f5",
    x"a1", x"fd", x"21", x"42", x"36", x"2e", x"32", x"06",
    x"10", x"e8", x"fc", x"31", x"b4", x"a2", x"0c", x"b7",
    x"b5", x"d0", x"ff", x"eb", x"0c", x"d8", x"f5", x"f7",
    x"f1", x"3d", x"2f", x"83", x"22", x"3b", x"cb", x"c0",
    x"fa", x"df", x"e1", x"93", x"ba", x"ee", x"d8", x"26",
    x"03", x"10", x"d4", x"c6", x"cc", x"a5", x"33", x"4e",
    x"ce", x"68", x"5f", x"ff", x"08", x"00", x"f9", x"09",
    x"01", x"fc", x"09", x"02", x"02", x"7a", x"b5", x"a9",
    x"96", x"b4", x"ab", x"fd", x"0c", x"3e", x"13", x"13",
    x"22", x"1d", x"25", x"06", x"ff", x"f0", x"ff", x"0c",
    x"02", x"f4", x"f8", x"10", x"f2", x"03", x"fe", x"c7",
    x"d0", x"dd", x"d9", x"fa", x"06", x"12", x"fc", x"f9",
    x"07", x"e9", x"c6", x"19", x"20", x"e1", x"13", x"fe",
    x"fe", x"c7", x"ad", x"df", x"01", x"31", x"30", x"f9",
    x"13", x"13", x"e7", x"11", x"2a", x"09", x"05", x"fa",
    x"27", x"14", x"e1", x"eb", x"0d", x"ef", x"10", x"34",
    x"1f", x"e8", x"50", x"2f", x"01", x"04", x"03", x"03",
    x"03", x"07", x"09", x"06", x"02", x"e4", x"f0", x"a8",
    x"f4", x"b1", x"ac", x"df", x"07", x"16", x"1e", x"b7",
    x"84", x"1c", x"ac", x"a2", x"d9", x"e4", x"f5", x"2a",
    x"14", x"0e", x"d8", x"b6", x"b2", x"d5", x"c5", x"0b",
    x"ff", x"fd", x"fe", x"ff", x"fd", x"02", x"fe", x"06",
    x"02", x"10", x"f6", x"df", x"a7", x"ca", x"d9", x"d4",
    x"f5", x"12", x"93", x"cc", x"e4", x"9f", x"10", x"01",
    x"16", x"1d", x"20", x"f5", x"ea", x"15", x"f6", x"2f",
    x"31", x"30", x"46", x"33", x"d8", x"c6", x"f2", x"ea",
    x"07", x"d4", x"fe", x"14", x"0d", x"e2", x"00", x"2a",
    x"1a", x"fd", x"0a", x"fb", x"20", x"1e", x"b3", x"d0",
    x"f5", x"64", x"05", x"0c", x"82", x"0c", x"19", x"2a",
    x"11", x"de", x"38", x"0c", x"18", x"16", x"14", x"e9",
    x"ff", x"fd", x"fb", x"fd", x"ff", x"fc", x"03", x"02",
    x"ff", x"01", x"fd", x"03", x"ff", x"00", x"04", x"fd",
    x"fe", x"04", x"42", x"29", x"19", x"09", x"09", x"08",
    x"30", x"0c", x"fc", x"d2", x"24", x"b0", x"25", x"22",
    x"e7", x"1b", x"1d", x"fe", x"2e", x"f7", x"e7", x"ef",
    x"ea", x"e8", x"ed", x"be", x"d6", x"c5", x"bc", x"04",
    x"f1", x"1a", x"1e", x"bd", x"2a", x"08", x"3a", x"23",
    x"25", x"cd", x"bf", x"cb", x"78", x"c0", x"d5", x"33",
    x"fe", x"2f", x"51", x"3c", x"0c", x"26", x"11", x"e8",
    x"31", x"16", x"30", x"1f", x"0c", x"c7", x"32", x"b2",
    x"c0", x"ed", x"e8", x"f4", x"ea", x"db", x"de", x"1d",
    x"ee", x"d3", x"f7", x"16", x"32", x"21", x"e4", x"ba",
    x"33", x"c1", x"d4", x"22", x"fc", x"d9", x"d7", x"eb",
    x"ca", x"d9", x"06", x"ff", x"0a", x"57", x"1f", x"30",
    x"32", x"39", x"33", x"16", x"1b", x"db", x"da", x"08",
    x"e6", x"f0", x"ea", x"18", x"11", x"ed", x"fa", x"2b",
    x"3e", x"d2", x"13", x"0e", x"01", x"fa", x"e4", x"7c",
    x"2b", x"fe", x"15", x"08", x"1e", x"f8", x"e7", x"f5",
    x"ef", x"2c", x"1f", x"e8", x"06", x"ec", x"d7", x"f3",
    x"53", x"e1", x"27", x"32", x"d8", x"df", x"e1", x"b8",
    x"f7", x"06", x"b2", x"d5", x"fc", x"fb", x"1d", x"1c",
    x"2f", x"28", x"21", x"fd", x"c2", x"e7", x"fb", x"14",
    x"d4", x"16", x"18", x"f1", x"d6", x"02", x"11", x"ac",
    x"0c", x"14", x"0f", x"24", x"3b", x"04", x"18", x"e6",
    x"c7", x"f2", x"f1", x"8c", x"e0", x"ee", x"e5", x"29",
    x"31", x"bc", x"d9", x"15", x"1f", x"ee", x"23", x"2d",
    x"0e", x"06", x"07", x"fa", x"01", x"06", x"02", x"f1",
    x"04", x"32", x"56", x"25", x"2b", x"3a", x"0c", x"0e",
    x"ec", x"01", x"1a", x"f6", x"1e", x"15", x"fb", x"c9",
    x"e0", x"d0", x"42", x"5f", x"20", x"0a", x"36", x"36",
    x"06", x"f5", x"0e", x"a2", x"b1", x"0e", x"9f", x"9e",
    x"f5", x"9d", x"e7", x"fa", x"40", x"0d", x"e7", x"ee",
    x"ff", x"ea", x"0c", x"f4", x"1d", x"2a", x"ff", x"37",
    x"fc", x"ec", x"e9", x"fe", x"e6", x"d8", x"95", x"a6",
    x"d3", x"a5", x"e9", x"0f", x"d9", x"f6", x"01", x"cf",
    x"00", x"90", x"47", x"4a", x"cd", x"49", x"f3", x"a7",
    x"34", x"39", x"18", x"05", x"12", x"e0", x"5b", x"d8",
    x"dd", x"01", x"06", x"04", x"02", x"04", x"05", x"fc",
    x"fe", x"00", x"44", x"ee", x"0d", x"c6", x"1c", x"07",
    x"12", x"fa", x"fb", x"0a", x"19", x"19", x"ef", x"e9",
    x"df", x"b3", x"e5", x"bb", x"cc", x"e3", x"20", x"21",
    x"23", x"09", x"24", x"f5", x"ec", x"f2", x"1f", x"02",
    x"0e", x"3f", x"1e", x"3c", x"1b", x"04", x"2f", x"16",
    x"09", x"23", x"25", x"04", x"3d", x"50", x"63", x"d0",
    x"22", x"58", x"cc", x"10", x"35", x"4d", x"4c", x"49",
    x"26", x"ab", x"14", x"0b", x"7c", x"f9", x"2d", x"38",
    x"1f", x"b8", x"ca", x"1b", x"d0", x"e9", x"0e", x"8d",
    x"c5", x"d2", x"03", x"04", x"24", x"1d", x"02", x"fe",
    x"c3", x"cd", x"ff", x"04", x"fd", x"00", x"03", x"ff",
    x"fc", x"04", x"0b", x"ff", x"41", x"53", x"16", x"23",
    x"0d", x"27", x"f6", x"fc", x"ee", x"11", x"16", x"11",
    x"a5", x"e8", x"f2", x"f4", x"fc", x"e8", x"d2", x"cd",
    x"e8", x"24", x"f8", x"e9", x"f5", x"18", x"0a", x"df",
    x"1a", x"21", x"0a", x"21", x"15", x"df", x"17", x"e2",
    x"d3", x"0e", x"2e", x"f3", x"bc", x"13", x"a4", x"c0",
    x"65", x"0b", x"15", x"29", x"fc", x"05", x"22", x"d6",
    x"c1", x"cf", x"ea", x"df", x"ba", x"b7", x"98", x"74",
    x"98", x"cb", x"f8", x"d1", x"24", x"f0", x"f9", x"04",
    x"f7", x"de", x"b6", x"c7", x"02", x"0c", x"07", x"04",
    x"00", x"03", x"fd", x"04", x"04", x"26", x"00", x"42",
    x"f5", x"f7", x"0a", x"fc", x"ff", x"d4", x"0a", x"97",
    x"f6", x"ff", x"fb", x"2f", x"3b", x"48", x"4e", x"2c",
    x"0b", x"52", x"bb", x"db", x"f7", x"8d", x"1d", x"11",
    x"fb", x"fe", x"03", x"00", x"00", x"00", x"05", x"03",
    x"03", x"07", x"b4", x"fa", x"b2", x"ea", x"04", x"ef",
    x"ba", x"b9", x"06", x"fa", x"1d", x"04", x"f4", x"1d",
    x"fc", x"0c", x"31", x"ed", x"18", x"e4", x"d9", x"d7",
    x"e1", x"37", x"f7", x"ea", x"15", x"0b", x"27", x"84",
    x"22", x"21", x"fd", x"2e", x"0a", x"d3", x"05", x"32",
    x"14", x"33", x"2f", x"f9", x"20", x"fa", x"45", x"f7",
    x"d0", x"e9", x"ab", x"d8", x"f8", x"d8", x"c2", x"d5",
    x"f1", x"11", x"02", x"07", x"03", x"15", x"fc", x"ee",
    x"06", x"03", x"fd", x"04", x"ff", x"04", x"06", x"01",
    x"00", x"fc", x"fa", x"04", x"ff", x"fd", x"02", x"fe",
    x"08", x"fa", x"04", x"f1", x"d2", x"01", x"f5", x"0f",
    x"09", x"17", x"27", x"16", x"d1", x"36", x"c7", x"06",
    x"3d", x"c6", x"02", x"4d", x"b7", x"0a", x"0f", x"79",
    x"c7", x"f9", x"af", x"d6", x"b9", x"f9", x"ed", x"02",
    x"c1", x"eb", x"f3", x"2e", x"f7", x"ce", x"14", x"ef",
    x"2f", x"36", x"da", x"12", x"d5", x"f3", x"08", x"14",
    x"d1", x"d9", x"ef", x"fa", x"1a", x"02", x"08", x"2f",
    x"e2", x"b2", x"08", x"bf", x"7c", x"ef", x"aa", x"c6",
    x"36", x"51", x"fd", x"04", x"ca", x"c4", x"d8", x"a4",
    x"b2", x"ff", x"ff", x"a3", x"b2", x"01", x"ed", x"e4",
    x"10", x"ee", x"00", x"0d", x"2f", x"fc", x"cd", x"ec",
    x"11", x"a1", x"ae", x"e6", x"22", x"fd", x"f5", x"d3",
    x"ff", x"dc", x"dd", x"e6", x"cd", x"0f", x"2b", x"20",
    x"ff", x"d9", x"d4", x"00", x"c9", x"bc", x"03", x"d9",
    x"94", x"17", x"e2", x"e2", x"d9", x"07", x"fa", x"f0",
    x"fe", x"e5", x"22", x"f4", x"cb", x"0e", x"ed", x"16",
    x"12", x"0f", x"e5", x"1a", x"37", x"d2", x"3a", x"33",
    x"08", x"23", x"07", x"15", x"09", x"1a", x"f8", x"fe",
    x"f1", x"bf", x"2c", x"22", x"ff", x"fc", x"fa", x"fe",
    x"ba", x"d0", x"0a", x"c3", x"ec", x"07", x"b1", x"cd",
    x"e8", x"e7", x"fc", x"d0", x"da", x"ec", x"ff", x"c9",
    x"d9", x"f8", x"83", x"c2", x"e2", x"f7", x"00", x"fb",
    x"19", x"21", x"35", x"05", x"26", x"3c", x"20", x"09",
    x"06", x"36", x"e1", x"e1", x"71", x"57", x"9f", x"5c",
    x"aa", x"e3", x"f1", x"0c", x"5d", x"3a", x"3f", x"32",
    x"c7", x"c5", x"b2", x"05", x"06", x"4a", x"10", x"08",
    x"35", x"1e", x"02", x"f3", x"b0", x"c8", x"da", x"ab",
    x"01", x"ff", x"21", x"6c", x"2b", x"f0", x"07", x"f5",
    x"1b", x"e3", x"92", x"2d", x"10", x"2c", x"39", x"e2",
    x"fb", x"5f", x"66", x"ba", x"04", x"fd", x"06", x"fd",
    x"e3", x"f6", x"04", x"ec", x"fd", x"dd", x"14", x"33",
    x"e9", x"04", x"15", x"eb", x"ee", x"e1", x"ce", x"d2",
    x"c1", x"b0", x"ae", x"f6", x"06", x"de", x"06", x"f9",
    x"df", x"d4", x"c3", x"e2", x"ed", x"e1", x"1f", x"02",
    x"f1", x"0d", x"e1", x"1c", x"ef", x"f8", x"ce", x"e5",
    x"d6", x"01", x"ff", x"fc", x"fe", x"fc", x"fe", x"fe",
    x"05", x"fe", x"81", x"f1", x"00", x"e4", x"15", x"28",
    x"26", x"14", x"11", x"e5", x"0a", x"00", x"e2", x"f5",
    x"20", x"eb", x"18", x"35", x"1f", x"4a", x"73", x"15",
    x"4c", x"23", x"43", x"26", x"2d", x"e2", x"fa", x"30",
    x"22", x"3e", x"57", x"ef", x"08", x"32", x"08", x"08",
    x"16", x"d0", x"c3", x"d4", x"e1", x"f3", x"0b", x"07",
    x"04", x"17", x"f6", x"de", x"15", x"05", x"c9", x"e1",
    x"1f", x"3a", x"24", x"38", x"db", x"f4", x"c9", x"89",
    x"ad", x"f6", x"25", x"19", x"20", x"28", x"14", x"1f",
    x"1c", x"c6", x"ef", x"fd", x"09", x"2d", x"51", x"44",
    x"f8", x"df", x"d6", x"02", x"fe", x"fb", x"fb", x"fe",
    x"fe", x"00", x"00", x"fd", x"01", x"e1", x"de", x"f1",
    x"05", x"fd", x"09", x"ea", x"fb", x"39", x"06", x"18",
    x"56", x"2c", x"38", x"bb", x"1f", x"0e", x"19", x"09",
    x"df", x"b8", x"a5", x"ad", x"c0", x"cb", x"f6", x"d3",
    x"d6", x"e0", x"f8", x"fe", x"10", x"2a", x"2c", x"20",
    x"fb", x"f3", x"21", x"14", x"09", x"95", x"06", x"e9",
    x"47", x"fb", x"d9", x"e4", x"f1", x"07", x"08", x"e2",
    x"e8", x"0c", x"30", x"27", x"2b", x"30", x"07", x"fb",
    x"45", x"12", x"1f", x"eb", x"35", x"02", x"19", x"2d",
    x"1d", x"2e", x"ff", x"fa", x"11", x"07", x"fa", x"03",
    x"07", x"0f", x"05", x"07", x"07", x"03", x"10", x"21",
    x"0d", x"15", x"12", x"e3", x"07", x"cf", x"21", x"c2",
    x"d9", x"0f", x"b9", x"e7", x"01", x"d3", x"d0", x"16",
    x"c2", x"e9", x"12", x"06", x"e0", x"01", x"87", x"54",
    x"ff", x"02", x"04", x"fd", x"fc", x"ff", x"00", x"fd",
    x"04", x"2d", x"fe", x"e7", x"15", x"33", x"ff", x"fa",
    x"18", x"2e", x"df", x"da", x"ea", x"f1", x"1a", x"16",
    x"0d", x"25", x"10", x"45", x"25", x"15", x"f7", x"da",
    x"c8", x"de", x"84", x"95", x"dc", x"39", x"29", x"f6",
    x"01", x"25", x"d2", x"e8", x"0f", x"15", x"40", x"2a",
    x"f1", x"ef", x"d8", x"d2", x"d8", x"ea", x"db", x"32",
    x"18", x"dc", x"f6", x"1a", x"e7", x"0e", x"39", x"20",
    x"1b", x"fe", x"0e", x"f8", x"11", x"f1", x"fb", x"ff",
    x"01", x"ff", x"04", x"fc", x"01", x"ff", x"03", x"f9",
    x"fa", x"04", x"fd", x"05", x"ff", x"fe", x"ff", x"ff",
    x"07", x"04", x"23", x"f9", x"d4", x"17", x"21", x"1a",
    x"ec", x"fc", x"13", x"27", x"30", x"12", x"27", x"a8",
    x"4d", x"23", x"7d", x"36", x"1f", x"0f", x"03", x"38",
    x"eb", x"f8", x"ef", x"f5", x"12", x"f8", x"f3", x"13",
    x"21", x"33", x"47", x"1e", x"4a", x"15", x"fc", x"ec",
    x"ed", x"d9", x"e6", x"06", x"23", x"f6", x"14", x"20",
    x"2f", x"30", x"54", x"1a", x"02", x"00", x"29", x"e7",
    x"12", x"f4", x"cf", x"f4", x"e6", x"d6", x"11", x"94",
    x"71", x"09", x"f3", x"11", x"4d", x"38", x"da", x"f8",
    x"01", x"89", x"f3", x"d9", x"e4", x"f2", x"1b", x"1b",
    x"f8", x"fd", x"fb", x"05", x"39", x"30", x"ff", x"e3",
    x"ee", x"0d", x"1b", x"30", x"f6", x"d9", x"ce", x"42",
    x"2d", x"1a", x"0c", x"2e", x"31", x"3a", x"13", x"15",
    x"2a", x"f6", x"f8", x"1f", x"df", x"c7", x"a0", x"c4",
    x"ba", x"0e", x"15", x"00", x"33", x"2b", x"d8", x"28",
    x"4a", x"15", x"03", x"e6", x"b2", x"06", x"d7", x"df",
    x"35", x"55", x"a9", x"f0", x"ff", x"db", x"23", x"26",
    x"42", x"1b", x"2b", x"3f", x"ec", x"20", x"f3", x"e1",
    x"12", x"ef", x"8a", x"6e", x"83", x"bf", x"ac", x"b2",
    x"4e", x"50", x"30", x"f6", x"a6", x"e2", x"03", x"e3",
    x"d4", x"d0", x"a8", x"ce", x"fc", x"0b", x"0a", x"f7",
    x"ef", x"cf", x"fb", x"f5", x"00", x"2d", x"03", x"0f",
    x"01", x"19", x"15", x"f6", x"19", x"49", x"b7", x"e5",
    x"ba", x"ef", x"f9", x"ec", x"11", x"2b", x"44", x"20",
    x"5e", x"4b", x"13", x"c5", x"dc", x"be", x"b1", x"ef",
    x"14", x"28", x"fb", x"10", x"ea", x"c1", x"d2", x"e2",
    x"b3", x"23", x"13", x"08", x"60", x"31", x"3d", x"41",
    x"1b", x"ef", x"f6", x"c6", x"d3", x"16", x"f5", x"39",
    x"3f", x"fd", x"15", x"be", x"ee", x"08", x"90", x"fd",
    x"1f", x"f5", x"36", x"4f", x"49", x"29", x"34", x"18",
    x"0e", x"12", x"1d", x"0d", x"0b", x"d4", x"fb", x"0d",
    x"ed", x"11", x"05", x"04", x"ef", x"09", x"3e", x"16",
    x"25", x"f0", x"fe", x"d0", x"dd", x"cc", x"f1", x"f6",
    x"bd", x"b3", x"ea", x"fc", x"ed", x"0c", x"f4", x"34",
    x"28", x"25", x"2e", x"13", x"31", x"3c", x"f0", x"1e",
    x"2c", x"fd", x"fb", x"fd", x"fc", x"05", x"fd", x"04",
    x"03", x"05", x"66", x"4f", x"71", x"e8", x"06", x"ed",
    x"a8", x"bd", x"ce", x"f8", x"09", x"31", x"2f", x"13",
    x"2c", x"5d", x"1d", x"0a", x"fb", x"f5", x"fb", x"eb",
    x"11", x"47", x"fa", x"19", x"15", x"00", x"16", x"16",
    x"38", x"33", x"0c", x"da", x"dc", x"cf", x"f7", x"3a",
    x"36", x"12", x"4d", x"47", x"d4", x"fe", x"0a", x"18",
    x"45", x"ff", x"dd", x"10", x"f1", x"c7", x"fd", x"e2",
    x"03", x"0e", x"e0", x"b3", x"f6", x"f1", x"fa", x"14",
    x"06", x"c3", x"be", x"10", x"05", x"0f", x"32", x"1d",
    x"fc", x"f3", x"14", x"f6", x"f4", x"00", x"ff", x"07",
    x"0d", x"fe", x"df", x"04", x"03", x"05", x"03", x"05",
    x"03", x"01", x"ff", x"ff", x"00", x"3c", x"51", x"ed",
    x"06", x"e9", x"d6", x"db", x"f5", x"ef", x"de", x"da",
    x"20", x"08", x"ef", x"23", x"0b", x"00", x"eb", x"ec",
    x"13", x"08", x"ff", x"f1", x"03", x"ed", x"e0", x"22",
    x"f7", x"22", x"dc", x"d8", x"e6", x"0b", x"fb", x"e9",
    x"1f", x"45", x"0b", x"18", x"10", x"fa", x"0a", x"fd",
    x"d6", x"06", x"f9", x"18", x"1e", x"fd", x"1a", x"1a",
    x"2b", x"12", x"f0", x"d0", x"d4", x"a2", x"d4", x"e6",
    x"07", x"ef", x"f3", x"62", x"7e", x"02", x"4f", x"01",
    x"ed", x"24", x"0c", x"f6", x"04", x"fe", x"fd", x"02",
    x"03", x"02", x"01", x"f5", x"f7", x"29", x"3c", x"30",
    x"00", x"4c", x"5f", x"0c", x"2b", x"46", x"17", x"f6",
    x"e5", x"46", x"ff", x"e5", x"2b", x"ed", x"db", x"04",
    x"f7", x"e7", x"11", x"05", x"ed", x"37", x"3b", x"29",
    x"05", x"fc", x"01", x"fb", x"fd", x"04", x"02", x"ff",
    x"fe", x"cc", x"a5", x"73", x"b9", x"ac", x"a5", x"21",
    x"1f", x"1e", x"0d", x"f0", x"de", x"01", x"dd", x"a8",
    x"09", x"b9", x"fa", x"e3", x"f0", x"f8", x"e0", x"e8",
    x"f1", x"30", x"eb", x"e9", x"06", x"e7", x"dd", x"d4",
    x"27", x"46", x"e3", x"24", x"2e", x"26", x"01", x"1e",
    x"00", x"ec", x"e9", x"09", x"e4", x"04", x"19", x"71",
    x"1f", x"c8", x"09", x"fc", x"af", x"e3", x"e7", x"2d",
    x"53", x"50", x"0f", x"24", x"0a", x"12", x"13", x"16",
    x"00", x"00", x"03", x"00", x"fe", x"03", x"01", x"05",
    x"00", x"09", x"03", x"01", x"ff", x"05", x"00", x"00",
    x"02", x"01", x"38", x"3a", x"42", x"11", x"0d", x"3b",
    x"eb", x"13", x"e2", x"20", x"3b", x"f6", x"10", x"28",
    x"2d", x"22", x"03", x"d5", x"09", x"12", x"1c", x"25",
    x"19", x"40", x"19", x"15", x"22", x"06", x"0f", x"0f",
    x"e6", x"e9", x"ec", x"06", x"ee", x"ef", x"46", x"43",
    x"4f", x"0b", x"64", x"57", x"db", x"2e", x"39", x"a9",
    x"0c", x"fa", x"f2", x"a4", x"e3", x"2f", x"fb", x"fb",
    x"dd", x"0f", x"1d", x"db", x"14", x"0b", x"fb", x"09",
    x"1a", x"e5", x"d9", x"07", x"fe", x"0d", x"11", x"12",
    x"04", x"11", x"d4", x"e2", x"d1", x"1f", x"f3", x"0e",
    x"2c", x"12", x"31", x"05", x"b3", x"dc", x"2e", x"fe",
    x"eb", x"22", x"12", x"f1", x"f7", x"2a", x"18", x"0b",
    x"19", x"fc", x"17", x"2a", x"1f", x"e6", x"0e", x"fa",
    x"ca", x"01", x"e1", x"08", x"17", x"f9", x"1d", x"ef",
    x"dc", x"0d", x"08", x"a6", x"d6", x"f2", x"e1", x"9b",
    x"a9", x"c4", x"c4", x"b6", x"f1", x"16", x"04", x"05",
    x"0e", x"c9", x"cb", x"06", x"d1", x"0b", x"1f", x"14",
    x"f7", x"ea", x"db", x"ec", x"34", x"03", x"ca", x"1c",
    x"d2", x"b3", x"4e", x"09", x"e5", x"c8", x"fe", x"02",
    x"f7", x"0b", x"24", x"0c", x"f5", x"ed", x"eb", x"c8",
    x"1e", x"0a", x"4a", x"0c", x"4e", x"06", x"0c", x"dd",
    x"f4", x"d6", x"1b", x"21", x"1a", x"2c", x"2d", x"eb",
    x"28", x"0f", x"c4", x"3a", x"30", x"1d", x"f0", x"f0",
    x"0c", x"26", x"19", x"0f", x"05", x"25", x"29", x"82",
    x"c3", x"0c", x"3c", x"41", x"0f", x"13", x"1a", x"11",
    x"2a", x"09", x"d1", x"34", x"14", x"fe", x"0b", x"f7",
    x"f9", x"27", x"20", x"1a", x"99", x"d9", x"fb", x"a9",
    x"f8", x"0d", x"03", x"34", x"39", x"e3", x"ee", x"34",
    x"53", x"e1", x"f9", x"b1", x"95", x"18", x"ce", x"e4",
    x"1f", x"ed", x"cd", x"06", x"39", x"d7", x"c4", x"03",
    x"fc", x"ed", x"18", x"03", x"08", x"51", x"68", x"a4",
    x"cd", x"bc", x"34", x"11", x"ec", x"26", x"17", x"5c",
    x"6a", x"c0", x"1e", x"27", x"1f", x"13", x"12", x"fa",
    x"fc", x"05", x"cf", x"39", x"fa", x"04", x"19", x"f5",
    x"13", x"1c", x"f4", x"31", x"18", x"fe", x"23", x"f8",
    x"f3", x"fe", x"fd", x"05", x"00", x"02", x"05", x"02",
    x"02", x"02", x"ee", x"11", x"02", x"d6", x"f2", x"14",
    x"24", x"0f", x"e4", x"05", x"e3", x"e4", x"06", x"06",
    x"f9", x"a1", x"bc", x"d0", x"87", x"d8", x"c3", x"1c",
    x"1a", x"13", x"ee", x"fd", x"ec", x"05", x"0f", x"1c",
    x"1f", x"f4", x"02", x"09", x"a6", x"ab", x"18", x"0c",
    x"e8", x"42", x"2d", x"1a", x"15", x"03", x"ff", x"de",
    x"86", x"0f", x"eb", x"de", x"04", x"bf", x"c1", x"1a",
    x"b6", x"fd", x"7f", x"3b", x"ac", x"e1", x"46", x"e4",
    x"eb", x"04", x"18", x"40", x"2d", x"2b", x"1d", x"30",
    x"ef", x"04", x"f3", x"0b", x"19", x"05", x"f6", x"f3",
    x"c1", x"bb", x"c4", x"fe", x"00", x"ff", x"06", x"04",
    x"f3", x"f8", x"fd", x"f9", x"fc", x"db", x"07", x"0a",
    x"f9", x"49", x"d9", x"e7", x"30", x"35", x"14", x"3c",
    x"2a", x"0d", x"4a", x"fe", x"36", x"3a", x"ec", x"f3",
    x"eb", x"d9", x"01", x"08", x"0a", x"02", x"01", x"fb",
    x"02", x"17", x"1c", x"20", x"24", x"2b", x"1f", x"23",
    x"d0", x"f8", x"e1", x"2f", x"12", x"3a", x"21", x"1b",
    x"32", x"de", x"d9", x"1f", x"b1", x"c5", x"ec", x"bc",
    x"ec", x"25", x"14", x"2d", x"e2", x"06", x"f2", x"0e",
    x"42", x"0e", x"c9", x"27", x"7d", x"da", x"03", x"c0",
    x"e1", x"2e", x"ee", x"f1", x"ff", x"03", x"01", x"f4",
    x"02", x"fe", x"04", x"fd", x"02", x"f2", x"1b", x"24",
    x"e7", x"fd", x"fa", x"e2", x"f5", x"f4", x"f6", x"ec",
    x"e8", x"1b", x"1b", x"19", x"21", x"67", x"40", x"c3",
    x"04", x"07", x"d3", x"05", x"29", x"14", x"6c", x"54",
    x"fc", x"ff", x"01", x"fd", x"fc", x"01", x"fd", x"00",
    x"01", x"08", x"f0", x"ff", x"d4", x"2f", x"13", x"cf",
    x"fb", x"f0", x"ef", x"b1", x"01", x"c4", x"ef", x"00",
    x"06", x"e9", x"d9", x"02", x"f4", x"f8", x"22", x"e4",
    x"e3", x"d7", x"b0", x"f5", x"fb", x"06", x"f9", x"c3",
    x"c0", x"f1", x"0f", x"d5", x"ee", x"d2", x"e3", x"d3",
    x"fd", x"14", x"f7", x"00", x"f4", x"f8", x"16", x"c2",
    x"c4", x"f7", x"06", x"eb", x"d4", x"f8", x"f9", x"e1",
    x"e6", x"02", x"a0", x"c9", x"f8", x"f4", x"e1", x"f8",
    x"fe", x"08", x"05", x"06", x"ff", x"0a", x"01", x"06",
    x"fe", x"fa", x"f9", x"fe", x"05", x"00", x"f7", x"ff",
    x"02", x"f8", x"58", x"3b", x"1d", x"04", x"01", x"f4",
    x"1f", x"13", x"30", x"c8", x"01", x"26", x"f4", x"15",
    x"55", x"1a", x"fd", x"1f", x"00", x"09", x"0e", x"00",
    x"01", x"13", x"38", x"08", x"f4", x"f4", x"f4", x"33",
    x"20", x"0d", x"0e", x"42", x"01", x"fe", x"c1", x"a5",
    x"f4", x"c5", x"c2", x"e6", x"30", x"e9", x"0a", x"f9",
    x"94", x"97", x"59", x"07", x"f0", x"4c", x"53", x"16",
    x"e8", x"1b", x"f4", x"1d", x"ea", x"1d", x"12", x"e8",
    x"0d", x"0a", x"13", x"18", x"0f", x"19", x"fb", x"fd",
    x"cb", x"c8", x"b6", x"0a", x"fb", x"03", x"11", x"18",
    x"03", x"17", x"27", x"fd", x"28", x"09", x"e9", x"0c",
    x"ed", x"0a", x"02", x"f0", x"0c", x"e3", x"b5", x"da",
    x"dc", x"f7", x"c9", x"ca", x"ff", x"15", x"03", x"f8",
    x"f8", x"ff", x"14", x"cf", x"d5", x"ff", x"07", x"1e",
    x"de", x"26", x"f2", x"ac", x"39", x"f6", x"dc", x"3b",
    x"0b", x"f0", x"28", x"29", x"14", x"1a", x"07", x"25",
    x"42", x"13", x"e0", x"13", x"1f", x"f4", x"15", x"31",
    x"1b", x"1b", x"25", x"0c", x"b3", x"1a", x"2e", x"ea",
    x"24", x"1f", x"09", x"fd", x"fd", x"1a", x"1c", x"21",
    x"28", x"f0", x"32", x"21", x"fe", x"19", x"05", x"03",
    x"16", x"13", x"3f", x"1d", x"e2", x"b3", x"0e", x"eb",
    x"e8", x"ce", x"d2", x"de", x"1b", x"19", x"e8", x"f4",
    x"15", x"08", x"c2", x"c4", x"c7", x"9a", x"a1", x"10",
    x"f8", x"69", x"ff", x"ec", x"f5", x"e5", x"0b", x"36",
    x"3e", x"d4", x"18", x"2b", x"ef", x"e4", x"fd", x"d6",
    x"19", x"f0", x"18", x"f9", x"0a", x"12", x"f8", x"f7",
    x"c1", x"f9", x"09", x"1e", x"08", x"bc", x"73", x"6a",
    x"38", x"af", x"13", x"0d", x"01", x"01", x"eb", x"e3",
    x"0a", x"13", x"f4", x"01", x"f7", x"e1", x"05", x"fd",
    x"0b", x"12", x"04", x"ff", x"09", x"ed", x"fb", x"0a",
    x"11", x"f1", x"30", x"de", x"e7", x"1b", x"16", x"61",
    x"18", x"0b", x"9d", x"ee", x"fd", x"d5", x"0d", x"fb",
    x"23", x"c6", x"e2", x"20", x"d6", x"b2", x"e7", x"0d",
    x"1c", x"dc", x"28", x"21", x"1f", x"3d", x"13", x"fb",
    x"d3", x"b3", x"fe", x"f5", x"24", x"0d", x"f5", x"d0",
    x"56", x"ff", x"ff", x"03", x"04", x"02", x"fe", x"fe",
    x"05", x"01", x"9e", x"b5", x"e4", x"b2", x"b4", x"cb",
    x"c9", x"b0", x"8b", x"02", x"1f", x"29", x"1f", x"f9",
    x"3b", x"d7", x"c5", x"f5", x"19", x"45", x"20", x"31",
    x"40", x"1c", x"2f", x"56", x"23", x"ec", x"01", x"fc",
    x"a2", x"c1", x"f9", x"76", x"64", x"9d", x"e8", x"d3",
    x"c4", x"da", x"f9", x"e6", x"cc", x"fd", x"00", x"fb",
    x"e6", x"fb", x"de", x"d3", x"fe", x"cc", x"c5", x"d5",
    x"e1", x"11", x"fc", x"ab", x"25", x"f3", x"cb", x"10",
    x"0c", x"0c", x"f9", x"25", x"d1", x"fc", x"0c", x"d3",
    x"31", x"50", x"19", x"ef", x"ea", x"ee", x"f9", x"e9",
    x"b4", x"c2", x"a3", x"0b", x"09", x"04", x"0b", x"01",
    x"05", x"07", x"fe", x"06", x"f1", x"eb", x"f5", x"f5",
    x"b0", x"a9", x"ef", x"d7", x"e5", x"f6", x"fa", x"30",
    x"02", x"ee", x"54", x"1a", x"41", x"37", x"13", x"10",
    x"ec", x"04", x"27", x"29", x"6d", x"30", x"27", x"da",
    x"be", x"e0", x"98", x"80", x"da", x"04", x"dd", x"9f",
    x"02", x"ff", x"fb", x"0e", x"22", x"fb", x"01", x"fa",
    x"fc", x"f9", x"07", x"27", x"e3", x"92", x"62", x"06",
    x"04", x"83", x"55", x"58", x"2b", x"ea", x"17", x"2a",
    x"ec", x"14", x"10", x"65", x"43", x"17", x"46", x"31",
    x"33", x"0e", x"1d", x"07", x"00", x"02", x"fe", x"fc",
    x"07", x"0b", x"fc", x"fc", x"fe", x"10", x"0d", x"d9",
    x"f8", x"0c", x"10", x"3c", x"01", x"04", x"01", x"2d",
    x"f8", x"f1", x"ff", x"ed", x"f4", x"0d", x"0c", x"d9",
    x"f0", x"ef", x"c6", x"dc", x"e0", x"db", x"03", x"f8",
    x"fb", x"fd", x"03", x"fd", x"00", x"02", x"00", x"fb",
    x"fb", x"47", x"37", x"0d", x"2f", x"4a", x"33", x"0e",
    x"22", x"40", x"c2", x"ea", x"cf", x"e9", x"d2", x"bb",
    x"07", x"d9", x"bd", x"13", x"19", x"19", x"d4", x"f1",
    x"ec", x"bd", x"46", x"1e", x"d5", x"db", x"a7", x"ca",
    x"ad", x"f5", x"ef", x"02", x"0e", x"1b", x"24", x"38",
    x"0a", x"2b", x"54", x"00", x"2c", x"2b", x"d8", x"fe",
    x"d1", x"a9", x"ef", x"f5", x"e1", x"d6", x"c5", x"b9",
    x"ab", x"e3", x"d0", x"d6", x"c1", x"a2", x"c9", x"bf",
    x"01", x"02", x"02", x"04", x"00", x"fd", x"fb", x"05",
    x"03", x"fe", x"03", x"03", x"01", x"01", x"fe", x"fd",
    x"03", x"01", x"02", x"1a", x"f3", x"d6", x"e7", x"ec",
    x"0f", x"d9", x"12", x"e5", x"06", x"77", x"f1", x"e4",
    x"db", x"ce", x"e9", x"cc", x"f6", x"f9", x"dd", x"15",
    x"f3", x"e0", x"fe", x"19", x"1c", x"be", x"b9", x"cc",
    x"cd", x"c8", x"e8", x"f0", x"7e", x"a3", x"22", x"f5",
    x"0c", x"dd", x"d7", x"c9", x"c1", x"0a", x"0d", x"13",
    x"14", x"fd", x"f3", x"07", x"14", x"19", x"00", x"12",
    x"de", x"14", x"ec", x"ea", x"e3", x"d5", x"e3", x"2d",
    x"14", x"bd", x"ca", x"f0", x"03", x"f0", x"f9", x"03",
    x"1a", x"2e", x"fb", x"b4", x"99", x"02", x"f4", x"1c",
    x"09", x"fa", x"f9", x"f3", x"e8", x"be", x"cf", x"ac",
    x"aa", x"f7", x"fa", x"be", x"08", x"f5", x"d6", x"22",
    x"eb", x"e2", x"66", x"21", x"26", x"fa", x"12", x"01",
    x"fe", x"24", x"0e", x"f0", x"fd", x"1b", x"34", x"43",
    x"fe", x"40", x"41", x"37", x"cc", x"37", x"12", x"2b",
    x"db", x"cf", x"e1", x"df", x"d3", x"0c", x"f4", x"a8",
    x"e2", x"16", x"cd", x"f5", x"11", x"ff", x"00", x"d8",
    x"fc", x"38", x"11", x"f5", x"df", x"e5", x"e8", x"e1",
    x"fe", x"07", x"f3", x"fa", x"1b", x"01", x"15", x"1b",
    x"06", x"1b", x"3e", x"09", x"fc", x"09", x"f9", x"28",
    x"06", x"e9", x"ee", x"d0", x"18", x"19", x"44", x"46",
    x"29", x"4c", x"21", x"59", x"53", x"86", x"0a", x"00",
    x"a8", x"d7", x"f1", x"1e", x"df", x"ed", x"c0", x"ce",
    x"e6", x"fb", x"ec", x"0f", x"00", x"2b", x"1c", x"3e",
    x"40", x"0c", x"35", x"29", x"06", x"24", x"10", x"e1",
    x"22", x"23", x"1e", x"25", x"21", x"06", x"00", x"05",
    x"cb", x"f6", x"df", x"ed", x"d8", x"cb", x"ee", x"d2",
    x"eb", x"1c", x"c6", x"ff", x"38", x"dc", x"45", x"54",
    x"10", x"1a", x"37", x"d3", x"d7", x"25", x"1d", x"f9",
    x"34", x"ec", x"14", x"21", x"15", x"fe", x"eb", x"0a",
    x"fb", x"f4", x"2d", x"0e", x"12", x"cf", x"e0", x"10",
    x"f3", x"ea", x"ce", x"fd", x"03", x"0c", x"23", x"5f",
    x"0f", x"15", x"22", x"1c", x"30", x"26", x"ee", x"33",
    x"1f", x"f3", x"30", x"22", x"e4", x"40", x"21", x"0d",
    x"23", x"e3", x"d7", x"25", x"db", x"e1", x"1f", x"ec",
    x"e0", x"fc", x"02", x"fe", x"fb", x"fc", x"fc", x"04",
    x"03", x"05", x"9a", x"fc", x"38", x"ff", x"30", x"25",
    x"13", x"01", x"f4", x"c4", x"e9", x"03", x"e0", x"f1",
    x"cf", x"bc", x"b7", x"c2", x"cf", x"bb", x"ce", x"1e",
    x"fc", x"fc", x"0c", x"ee", x"e7", x"f0", x"d7", x"fd",
    x"f0", x"db", x"d9", x"13", x"fe", x"e3", x"dd", x"e6",
    x"e3", x"1b", x"13", x"f9", x"41", x"26", x"13", x"22",
    x"3d", x"40", x"1a", x"2f", x"34", x"ed", x"13", x"4b",
    x"16", x"d6", x"e1", x"07", x"21", x"10", x"05", x"0f",
    x"1d", x"f7", x"e7", x"0d", x"d1", x"d5", x"df", x"a4",
    x"ce", x"f6", x"ff", x"f5", x"fa", x"e3", x"e4", x"cc",
    x"d3", x"e4", x"d1", x"01", x"08", x"00", x"fb", x"08",
    x"06", x"ff", x"05", x"f7", x"57", x"6a", x"7b", x"31",
    x"2d", x"52", x"23", x"45", x"3f", x"f8", x"1f", x"f2",
    x"f0", x"14", x"11", x"e8", x"e8", x"ca", x"18", x"cc",
    x"f1", x"21", x"23", x"1e", x"35", x"15", x"1c", x"3e",
    x"4e", x"40", x"2e", x"3a", x"4c", x"1b", x"f8", x"06",
    x"09", x"05", x"0d", x"a6", x"c5", x"ff", x"fa", x"01",
    x"57", x"d9", x"e8", x"0b", x"b9", x"cf", x"03", x"00",
    x"ea", x"cd", x"a8", x"d9", x"f9", x"dd", x"ed", x"18",
    x"d7", x"f2", x"fe", x"e1", x"05", x"17", x"15", x"c0",
    x"cc", x"e9", x"ba", x"c1", x"0e", x"09", x"08", x"0f",
    x"07", x"0f", x"0d", x"1c", x"0b", x"fb", x"f0", x"ec",
    x"0a", x"ce", x"be", x"2d", x"c8", x"c4", x"10", x"3c",
    x"49", x"10", x"50", x"25", x"25", x"2d", x"28", x"aa",
    x"e3", x"d9", x"0d", x"1f", x"1f", x"14", x"1f", x"26",
    x"02", x"fc", x"fc", x"fc", x"fd", x"fe", x"04", x"ff",
    x"fd", x"e2", x"f9", x"24", x"eb", x"fe", x"fe", x"24",
    x"cc", x"b4", x"e0", x"1a", x"41", x"fc", x"f9", x"1c",
    x"10", x"00", x"11", x"1a", x"28", x"17", x"0d", x"08",
    x"0b", x"d6", x"eb", x"09", x"44", x"16", x"0b", x"dd",
    x"af", x"a8", x"e6", x"c0", x"be", x"f8", x"f4", x"fa",
    x"e7", x"f9", x"ed", x"ef", x"c4", x"d9", x"f8", x"ae",
    x"fe", x"23", x"fa", x"fd", x"ff", x"d5", x"d4", x"84",
    x"61", x"c0", x"9e", x"a2", x"db", x"df", x"19", x"17",
    x"00", x"fe", x"ff", x"08", x"fc", x"05", x"fb", x"fb",
    x"05", x"00", x"fc", x"00", x"ff", x"02", x"fd", x"f8",
    x"00", x"fb", x"ea", x"01", x"f3", x"1c", x"1b", x"04",
    x"08", x"03", x"d0", x"a1", x"87", x"bc", x"cd", x"01",
    x"0c", x"dc", x"04", x"2a", x"90", x"a4", x"96", x"b9",
    x"6c", x"93", x"08", x"18", x"07", x"06", x"11", x"1f",
    x"13", x"1c", x"09", x"f4", x"f8", x"00", x"db", x"04",
    x"f1", x"bb", x"e4", x"d0", x"0d", x"f9", x"d5", x"97",
    x"75", x"92", x"f1", x"e4", x"ef", x"14", x"14", x"23",
    x"fd", x"cd", x"16", x"fe", x"f6", x"2c", x"d4", x"20",
    x"2f", x"fd", x"eb", x"06", x"92", x"c2", x"ef", x"a2",
    x"e2", x"03", x"d2", x"ad", x"dc", x"f5", x"08", x"05",
    x"c3", x"12", x"17", x"dc", x"e0", x"df", x"14", x"16",
    x"14", x"fd", x"25", x"30", x"09", x"09", x"21", x"d3",
    x"ac", x"f2", x"d1", x"cc", x"da", x"05", x"1b", x"31",
    x"ec", x"07", x"00", x"33", x"05", x"09", x"16", x"02",
    x"09", x"05", x"eb", x"f5", x"11", x"fb", x"05", x"c5",
    x"9f", x"ea", x"06", x"e1", x"dd", x"ff", x"08", x"0e",
    x"3e", x"23", x"2c", x"e0", x"eb", x"1e", x"e8", x"ff",
    x"2e", x"c5", x"e9", x"fa", x"a4", x"de", x"11", x"c6",
    x"db", x"ea", x"2f", x"10", x"49", x"20", x"0d", x"13",
    x"32", x"23", x"05", x"e0", x"c2", x"ec", x"fd", x"fb",
    x"24", x"fe", x"e7", x"de", x"d7", x"f8", x"0c", x"e8",
    x"b4", x"8e", x"03", x"ff", x"e1", x"17", x"fa", x"17",
    x"2d", x"36", x"3c", x"b8", x"36", x"1c", x"2a", x"e1",
    x"d5", x"27", x"3a", x"26", x"52", x"38", x"29", x"1e",
    x"1c", x"17", x"24", x"f3", x"c6", x"92", x"93", x"c8",
    x"1a", x"fd", x"ff", x"0b", x"e9", x"cd", x"d3", x"d0",
    x"cc", x"17", x"05", x"32", x"08", x"ee", x"ad", x"cf",
    x"0d", x"25", x"f4", x"e3", x"07", x"23", x"08", x"05",
    x"ff", x"2b", x"fb", x"36", x"03", x"01", x"00", x"41",
    x"30", x"17", x"52", x"24", x"20", x"0a", x"fc", x"0b",
    x"0a", x"13", x"47", x"1a", x"2a", x"15", x"f1", x"16",
    x"1d", x"0d", x"cf", x"1a", x"19", x"e7", x"fc", x"d6",
    x"13", x"58", x"3e", x"3b", x"5c", x"0d", x"18", x"28",
    x"0b", x"25", x"15", x"01", x"cb", x"28", x"0f", x"f3",
    x"06", x"2f", x"49", x"e0", x"03", x"14", x"c6", x"b1",
    x"c4", x"00", x"02", x"fd", x"ff", x"02", x"00", x"01",
    x"ff", x"fe", x"24", x"29", x"1a", x"09", x"ee", x"07",
    x"e1", x"ea", x"ee", x"f2", x"0c", x"ff", x"1f", x"16",
    x"f8", x"23", x"19", x"e8", x"e7", x"d7", x"ea", x"ef",
    x"f9", x"e9", x"82", x"d7", x"ef", x"0b", x"f8", x"09",
    x"f5", x"b6", x"d1", x"d9", x"f5", x"c3", x"08", x"1d",
    x"07", x"ef", x"fc", x"13", x"c9", x"ff", x"0a", x"20",
    x"e2", x"c9", x"08", x"a9", x"a9", x"b7", x"a7", x"c1",
    x"17", x"09", x"16", x"0b", x"f7", x"0d", x"ef", x"3a",
    x"1f", x"fe", x"e3", x"0b", x"eb", x"fe", x"e5", x"e1",
    x"eb", x"15", x"f4", x"f3", x"07", x"f1", x"ff", x"f1",
    x"f7", x"17", x"dd", x"05", x"f9", x"fe", x"08", x"fa",
    x"fb", x"00", x"ff", x"ff", x"1d", x"04", x"05", x"de",
    x"e9", x"d6", x"d0", x"d4", x"df", x"0d", x"e0", x"26",
    x"b8", x"ea", x"12", x"d6", x"e1", x"23", x"06", x"07",
    x"fa", x"5d", x"59", x"37", x"4c", x"da", x"d0", x"18",
    x"fb", x"09", x"13", x"f1", x"e3", x"a7", x"a8", x"26",
    x"e7", x"1f", x"e6", x"e2", x"27", x"23", x"fe", x"28",
    x"40", x"f6", x"0f", x"47", x"02", x"25", x"ec", x"18",
    x"0a", x"de", x"f5", x"f5", x"e6", x"0d", x"fc", x"e0",
    x"f9", x"fc", x"07", x"31", x"0a", x"e5", x"e9", x"cb",
    x"cd", x"ac", x"cb", x"ce", x"fd", x"01", x"fb", x"02",
    x"ff", x"02", x"01", x"f8", x"08", x"f0", x"f7", x"fb",
    x"df", x"ec", x"fd", x"df", x"f3", x"11", x"e5", x"01",
    x"1e", x"dc", x"18", x"19", x"5c", x"22", x"0c", x"e6",
    x"11", x"10", x"23", x"2e", x"4c", x"6f", x"37", x"3d",
    x"04", x"fc", x"fc", x"ff", x"01", x"04", x"fb", x"fe",
    x"03", x"1f", x"09", x"21", x"1e", x"04", x"02", x"0c",
    x"03", x"fd", x"1b", x"f5", x"11", x"ff", x"29", x"19",
    x"fb", x"18", x"04", x"3e", x"e2", x"e8", x"21", x"e7",
    x"d2", x"fd", x"99", x"a9", x"fc", x"f2", x"02", x"f2",
    x"df", x"ea", x"ed", x"d9", x"cb", x"fe", x"f4", x"f2",
    x"fd", x"e8", x"f2", x"ba", x"d8", x"e0", x"ee", x"08",
    x"1c", x"e1", x"7a", x"b3", x"05", x"e7", x"e7", x"17",
    x"f8", x"18", x"07", x"e2", x"12", x"02", x"05", x"05",
    x"fe", x"f5", x"fc", x"02", x"06", x"ff", x"ff", x"fc",
    x"ff", x"fa", x"f8", x"f9", x"01", x"00", x"02", x"02",
    x"04", x"f9", x"12", x"08", x"2b", x"d4", x"eb", x"ed",
    x"08", x"26", x"14", x"02", x"43", x"e2", x"1d", x"41",
    x"4e", x"21", x"13", x"db", x"fd", x"10", x"12", x"17",
    x"1e", x"09", x"ee", x"f3", x"1b", x"19", x"1e", x"10",
    x"22", x"c3", x"b1", x"da", x"91", x"cf", x"39", x"1c",
    x"18", x"15", x"3e", x"2b", x"03", x"f2", x"cc", x"09",
    x"13", x"07", x"f1", x"14", x"25", x"78", x"42", x"47",
    x"2f", x"1a", x"1d", x"e8", x"12", x"03", x"4a", x"2c",
    x"14", x"11", x"17", x"ff", x"a7", x"a6", x"bc", x"f0",
    x"9d", x"6b", x"2d", x"26", x"41", x"26", x"08", x"08",
    x"23", x"f7", x"29", x"04", x"0b", x"0b", x"26", x"1e",
    x"04", x"cd", x"e9", x"e1", x"db", x"2b", x"39", x"01",
    x"c7", x"c3", x"dc", x"18", x"19", x"0b", x"1e", x"07",
    x"27", x"b0", x"96", x"0d", x"6b", x"69", x"11", x"1a",
    x"1c", x"06", x"09", x"21", x"d2", x"08", x"f5", x"03",
    x"2c", x"13", x"e4", x"1e", x"13", x"f1", x"de", x"c7",
    x"eb", x"19", x"31", x"de", x"e8", x"d1", x"ef", x"de",
    x"3b", x"42", x"26", x"0c", x"50", x"1f", x"0e", x"20",
    x"23", x"0b", x"0a", x"20", x"31", x"e7", x"01", x"00",
    x"19", x"11", x"32", x"ff", x"f9", x"30", x"d6", x"d4",
    x"20", x"c2", x"ab", x"e6", x"07", x"14", x"0c", x"23",
    x"2b", x"ff", x"09", x"f9", x"e6", x"29", x"fd", x"30",
    x"fe", x"17", x"2b", x"05", x"19", x"10", x"d7", x"96",
    x"d2", x"ef", x"04", x"e6", x"0e", x"2c", x"34", x"eb",
    x"15", x"10", x"1d", x"21", x"34", x"03", x"07", x"08",
    x"3e", x"17", x"66", x"27", x"10", x"21", x"04", x"2d",
    x"17", x"de", x"26", x"21", x"04", x"2b", x"29", x"0c",
    x"0d", x"46", x"26", x"f9", x"04", x"23", x"22", x"27",
    x"5b", x"2b", x"e2", x"9e", x"c5", x"ed", x"9e", x"ea",
    x"e3", x"bd", x"f2", x"01", x"db", x"96", x"a9", x"05",
    x"f0", x"e6", x"0d", x"f4", x"00", x"2b", x"21", x"31",
    x"14", x"1e", x"37", x"08", x"e5", x"18", x"d7", x"d4",
    x"e1", x"f4", x"e7", x"f6", x"ef", x"ef", x"01", x"e1",
    x"ec", x"cf", x"f2", x"17", x"1b", x"04", x"22", x"57",
    x"e8", x"ef", x"05", x"e5", x"fe", x"31", x"f0", x"18",
    x"2f", x"02", x"01", x"fd", x"fb", x"fe", x"fb", x"01",
    x"ff", x"ff", x"01", x"0e", x"06", x"0e", x"f2", x"0a",
    x"03", x"14", x"09", x"22", x"51", x"59", x"0f", x"08",
    x"1b", x"20", x"0e", x"05", x"e4", x"3c", x"16", x"ff",
    x"3a", x"78", x"e3", x"1e", x"2d", x"26", x"e0", x"dd",
    x"44", x"ef", x"da", x"1f", x"f3", x"e9", x"16", x"e0",
    x"04", x"16", x"fe", x"fd", x"3b", x"f9", x"dd", x"15",
    x"07", x"ec", x"13", x"fd", x"26", x"03", x"f2", x"dd",
    x"04", x"d9", x"da", x"60", x"0b", x"fb", x"8d", x"0e",
    x"fa", x"03", x"0a", x"39", x"e9", x"13", x"14", x"17",
    x"1e", x"fb", x"51", x"28", x"2e", x"44", x"ed", x"00",
    x"09", x"bf", x"f7", x"0a", x"fb", x"fe", x"03", x"03",
    x"03", x"fa", x"fe", x"03", x"2a", x"f6", x"b3", x"29",
    x"f7", x"da", x"09", x"f5", x"f1", x"e1", x"c5", x"82",
    x"07", x"02", x"30", x"fa", x"ea", x"17", x"0a", x"f1",
    x"12", x"0b", x"18", x"1b", x"fb", x"1e", x"2b", x"f5",
    x"fb", x"d8", x"fd", x"fe", x"02", x"07", x"0f", x"11",
    x"a5", x"b2", x"f1", x"d0", x"da", x"84", x"d9", x"d8",
    x"95", x"13", x"1b", x"34", x"06", x"05", x"2c", x"e6",
    x"db", x"15", x"be", x"d8", x"06", x"ba", x"ce", x"d4",
    x"e4", x"ec", x"d9", x"12", x"3e", x"58", x"ed", x"10",
    x"22", x"26", x"14", x"0f", x"fe", x"fc", x"fc", x"05",
    x"02", x"fe", x"03", x"f9", x"02", x"5f", x"8e", x"84",
    x"16", x"60", x"56", x"2e", x"47", x"46", x"1a", x"1d",
    x"f3", x"ec", x"0f", x"ff", x"35", x"fb", x"f5", x"f3",
    x"e0", x"bb", x"17", x"c4", x"cb", x"0b", x"e6", x"f7",
    x"04", x"04", x"fb", x"fb", x"01", x"01", x"ff", x"04",
    x"01", x"15", x"56", x"23", x"39", x"33", x"1d", x"01",
    x"2c", x"20", x"42", x"73", x"61", x"2c", x"21", x"15",
    x"1d", x"ed", x"f8", x"42", x"19", x"01", x"53", x"1c",
    x"13", x"1e", x"12", x"08", x"49", x"44", x"3f", x"fb",
    x"2e", x"50", x"e6", x"17", x"34", x"0e", x"cb", x"ee",
    x"4f", x"27", x"16", x"29", x"36", x"e3", x"00", x"b3",
    x"89", x"ec", x"15", x"38", x"e8", x"ed", x"fd", x"30",
    x"ed", x"1e", x"0c", x"ec", x"fe", x"14", x"ee", x"f7",
    x"03", x"ff", x"fd", x"fe", x"fe", x"04", x"ff", x"00",
    x"01", x"06", x"05", x"ff", x"03", x"fe", x"fb", x"05",
    x"09", x"03", x"e5", x"9f", x"d8", x"e2", x"bd", x"f3",
    x"be", x"d3", x"e6", x"f9", x"7f", x"a1", x"ee", x"f7",
    x"d0", x"d6", x"f0", x"d0", x"21", x"06", x"e4", x"f9",
    x"df", x"f1", x"e5", x"e7", x"19", x"ef", x"e2", x"f9",
    x"e3", x"cc", x"f3", x"f2", x"96", x"bb", x"4a", x"c0",
    x"f1", x"e8", x"e6", x"fa", x"07", x"ff", x"00", x"b8",
    x"65", x"78", x"e0", x"f6", x"d4", x"0c", x"0c", x"0a",
    x"97", x"01", x"02", x"e3", x"03", x"fa", x"d1", x"37",
    x"15", x"e0", x"2a", x"f1", x"f6", x"06", x"ef", x"04",
    x"0f", x"05", x"13", x"04", x"e7", x"20", x"0a", x"e0",
    x"f4", x"17", x"00", x"07", x"10", x"12", x"0b", x"1d",
    x"ff", x"ef", x"17", x"03", x"4f", x"e3", x"04", x"15",
    x"10", x"1c", x"23", x"09", x"ff", x"0e", x"fb", x"ea",
    x"d7", x"fe", x"27", x"04", x"03", x"25", x"37", x"cb",
    x"ef", x"ff", x"15", x"02", x"e7", x"08", x"fc", x"d5",
    x"be", x"af", x"be", x"b6", x"96", x"05", x"e8", x"92",
    x"fa", x"fb", x"04", x"04", x"03", x"05", x"03", x"f9",
    x"ff", x"f7", x"03", x"fc", x"fd", x"00", x"03", x"fc",
    x"f8", x"fa", x"fe", x"05", x"fa", x"fd", x"01", x"fc",
    x"fa", x"00", x"fa", x"fa", x"fa", x"fc", x"f7", x"fc",
    x"f6", x"f9", x"f8", x"f3", x"01", x"02", x"ff", x"f8",
    x"00", x"ff", x"fd", x"fb", x"01", x"fb", x"f9", x"00",
    x"ff", x"fe", x"01", x"00", x"f7", x"fc", x"02", x"fc",
    x"03", x"f8", x"03", x"04", x"01", x"fc", x"01", x"04",
    x"fe", x"fe", x"fd", x"fc", x"fe", x"00", x"01", x"fb",
    x"03", x"02", x"ff", x"fc", x"ff", x"01", x"fe", x"fc",
    x"fb", x"00", x"00", x"fc", x"01", x"ff", x"02", x"fc",
    x"f7", x"fd", x"fc", x"ff", x"fa", x"01", x"fc", x"fc",
    x"00", x"f7", x"02", x"fd", x"fa", x"f9", x"f9", x"02",
    x"00", x"02", x"fe", x"01", x"f8", x"fe", x"01", x"fe",
    x"fd", x"03", x"fd", x"f9", x"fa", x"fd", x"fa", x"00",
    x"ff", x"02", x"fc", x"fc", x"01", x"04", x"fd", x"00",
    x"00", x"ff", x"fe", x"fe", x"00", x"fc", x"fe", x"fe",
    x"03", x"fa", x"fc", x"fe", x"fd", x"02", x"02", x"01",
    x"fd", x"fd", x"fe", x"fb", x"fd", x"fb", x"fb", x"03",
    x"fd", x"00", x"02", x"fd", x"fe", x"03", x"02", x"fe",
    x"04", x"fc", x"01", x"fa", x"fa", x"fd", x"ff", x"03",
    x"ff", x"01", x"01", x"f9", x"fc", x"fa", x"03", x"f8",
    x"fa", x"fa", x"fe", x"f8", x"f8", x"02", x"06", x"fc",
    x"00", x"fd", x"fe", x"00", x"fe", x"fc", x"fc", x"00",
    x"f9", x"03", x"ff", x"fc", x"f8", x"f9", x"fb", x"03",
    x"ff", x"fa", x"00", x"fe", x"03", x"fe", x"00", x"fe",
    x"ff", x"04", x"fb", x"fb", x"fd", x"00", x"fd", x"01",
    x"ff", x"f7", x"fe", x"fc", x"00", x"fc", x"f7", x"fd",
    x"ff", x"f7", x"fd", x"fc", x"fe", x"fc", x"04", x"fb",
    x"fc", x"fe", x"fd", x"f8", x"fd", x"02", x"fa", x"fc",
    x"ff", x"f4", x"02", x"00", x"00", x"03", x"00", x"ff",
    x"fd", x"04", x"00", x"fd", x"02", x"fb", x"03", x"fa",
    x"04", x"fb", x"00", x"02", x"ff", x"f9", x"02", x"04",
    x"fd", x"fd", x"04", x"fc", x"ff", x"04", x"fb", x"01",
    x"fd", x"fd", x"04", x"03", x"fd", x"ff", x"ff", x"03",
    x"04", x"fa", x"fa", x"00", x"fb", x"f7", x"fa", x"fd",
    x"03", x"fe", x"02", x"02", x"00", x"fc", x"fd", x"01",
    x"00", x"fb", x"fc", x"01", x"f5", x"fc", x"f6", x"fd",
    x"f5", x"fa", x"02", x"ff", x"00", x"01", x"01", x"fa",
    x"fe", x"03", x"fd", x"fc", x"f5", x"03", x"03", x"fd",
    x"fa", x"ff", x"fa", x"f8", x"06", x"05", x"02", x"00",
    x"fc", x"00", x"03", x"fb", x"00", x"03", x"04", x"03",
    x"fb", x"fa", x"02", x"ff", x"00", x"04", x"03", x"01",
    x"fa", x"fa", x"fc", x"01", x"01", x"f9", x"fe", x"fb",
    x"fc", x"fb", x"fb", x"03", x"fc", x"fa", x"fb", x"f9",
    x"fc", x"01", x"03", x"fd", x"02", x"04", x"ff", x"fe",
    x"06", x"fb", x"fe", x"fe", x"fb", x"01", x"04", x"fa",
    x"fd", x"fe", x"fd", x"fe", x"03", x"04", x"03", x"fd",
    x"03", x"fc", x"01", x"00", x"01", x"ff", x"05", x"f9",
    x"ff", x"fe", x"fc", x"03", x"fb", x"fa", x"fc", x"fd",
    x"04", x"fc", x"02", x"fa", x"fe", x"fb", x"02", x"02",
    x"01", x"fc", x"fa", x"fb", x"fc", x"fb", x"fe", x"04",
    x"fe", x"02", x"fc", x"ff", x"fc", x"03", x"fc", x"fd",
    x"fc", x"fc", x"fb", x"fb", x"01", x"04", x"fe", x"fa",
    x"fc", x"fd", x"fd", x"ff", x"fd", x"fd", x"ff", x"02",
    x"fc", x"05", x"fc", x"fb", x"fe", x"fc", x"02", x"01",
    x"fe", x"fd", x"fe", x"fe", x"02", x"ff", x"fc", x"fe",
    x"fd", x"02", x"fe", x"03", x"00", x"01", x"00", x"01",
    x"fc", x"fb", x"fb", x"fe", x"fa", x"05", x"fb", x"ff",
    x"fb", x"01", x"ff", x"fc", x"01", x"f9", x"fd", x"fa",
    x"f6", x"fd", x"03", x"f7", x"ff", x"fd", x"00", x"fd",
    x"fa", x"00", x"fa", x"fd", x"03", x"01", x"fe", x"fd",
    x"ff", x"ff", x"00", x"fe", x"00", x"02", x"f7", x"ff",
    x"fe", x"f6", x"ff", x"00", x"fb", x"fb", x"01", x"fd",
    x"ff", x"fe", x"ff", x"00", x"fa", x"fa", x"fe", x"05",
    x"00", x"fb", x"fa", x"f9", x"01", x"fe", x"fd", x"00",
    x"fa", x"f8", x"fd", x"f8", x"f9", x"fe", x"fd", x"fd",
    x"ff", x"fe", x"fd", x"fa", x"fc", x"00", x"00", x"fd",
    x"f7", x"fe", x"00", x"fb", x"ff", x"f7", x"fd", x"fd",
    x"fb", x"ff", x"fd", x"03", x"fb", x"01", x"fe", x"02",
    x"fe", x"fa", x"fb", x"01", x"01", x"00", x"01", x"f8",
    x"02", x"01", x"fd", x"fb", x"fb", x"f7", x"01", x"fe",
    x"3e", x"29", x"f8", x"4c", x"5a", x"21", x"15", x"22",
    x"05", x"0a", x"15", x"0b", x"ee", x"01", x"0e", x"bc",
    x"f3", x"b8", x"b4", x"dd", x"e9", x"dc", x"fc", x"fd",
    x"12", x"e5", x"02", x"07", x"1c", x"f2", x"24", x"19",
    x"fd", x"27", x"02", x"e8", x"fb", x"db", x"be", x"e3",
    x"b1", x"bc", x"b6", x"ff", x"e2", x"23", x"1e", x"20",
    x"30", x"07", x"b7", x"99", x"9e", x"c2", x"40", x"22",
    x"35", x"03", x"10", x"22", x"12", x"f7", x"00", x"41",
    x"35", x"57", x"d7", x"f8", x"0e", x"a8", x"d6", x"f5",
    x"f2", x"cc", x"bc", x"e1", x"e8", x"9a", x"fc", x"d9",
    x"e4", x"00", x"24", x"37", x"0c", x"16", x"27", x"ec",
    x"b0", x"81", x"31", x"f9", x"d4", x"50", x"2d", x"ec",
    x"f7", x"55", x"0f", x"18", x"f2", x"e9", x"c8", x"fc",
    x"e6", x"ff", x"e4", x"f0", x"df", x"2f", x"1d", x"e3",
    x"0e", x"fa", x"09", x"e2", x"04", x"e0", x"c0", x"e9",
    x"f2", x"d7", x"0b", x"df", x"f7", x"df", x"49", x"2a",
    x"47", x"ef", x"e2", x"ec", x"d8", x"e9", x"0f", x"de",
    x"a4", x"f0", x"db", x"d7", x"c1", x"f0", x"db", x"dd",
    x"d0", x"d2", x"ff", x"e1", x"e8", x"03", x"fc", x"fd",
    x"fd", x"01", x"fb", x"04", x"04", x"05", x"02", x"00",
    x"fc", x"fb", x"f6", x"00", x"cc", x"f5", x"ed", x"e7",
    x"e5", x"e3", x"f3", x"0a", x"29", x"0f", x"09", x"25",
    x"00", x"9a", x"16", x"5f", x"46", x"04", x"f0", x"10",
    x"fc", x"f6", x"84", x"ca", x"2f", x"fe", x"fa", x"0f",
    x"3e", x"2c", x"25", x"28", x"23", x"f9", x"fd", x"e5",
    x"d0", x"cc", x"09", x"eb", x"0e", x"18", x"31", x"07",
    x"a1", x"96", x"43", x"f4", x"ee", x"35", x"2c", x"0e",
    x"3f", x"e1", x"e5", x"e5", x"f8", x"eb", x"d1", x"ee",
    x"0f", x"1f", x"23", x"e4", x"34", x"2f", x"2c", x"be",
    x"fb", x"10", x"fa", x"02", x"23", x"22", x"33", x"34",
    x"be", x"b5", x"b7", x"06", x"03", x"07", x"03", x"02",
    x"05", x"fd", x"ff", x"fe", x"d3", x"bd", x"e0", x"f7",
    x"e7", x"14", x"10", x"f0", x"fc", x"be", x"20", x"57",
    x"1e", x"2e", x"0c", x"52", x"3b", x"37", x"d8", x"0f",
    x"0a", x"ae", x"c4", x"dc", x"ed", x"0d", x"d1", x"e4",
    x"09", x"e4", x"ab", x"c1", x"d8", x"8f", x"54", x"6a",
    x"7a", x"38", x"cf", x"50", x"16", x"ff", x"0c", x"f2",
    x"07", x"43", x"12", x"21", x"fe", x"f6", x"1b", x"e3",
    x"f9", x"fe", x"37", x"1e", x"2b", x"16", x"05", x"1b",
    x"81", x"f4", x"d9", x"49", x"3f", x"d8", x"34", x"20",
    x"1d", x"f6", x"ea", x"f1", x"f5", x"fd", x"00", x"f7",
    x"fc", x"05", x"f9", x"06", x"fe", x"d8", x"e0", x"b9",
    x"fc", x"1c", x"0b", x"1b", x"0c", x"0d", x"37", x"da",
    x"f4", x"19", x"eb", x"f6", x"f9", x"01", x"0e", x"db",
    x"15", x"15", x"fc", x"1a", x"1e", x"01", x"0a", x"1e",
    x"03", x"ff", x"04", x"fc", x"fc", x"fb", x"05", x"02",
    x"fd", x"9e", x"e1", x"f8", x"b3", x"e9", x"0d", x"f0",
    x"f5", x"1a", x"bf", x"89", x"ba", x"12", x"e4", x"f3",
    x"30", x"c5", x"c8", x"a5", x"e6", x"f1", x"01", x"24",
    x"e7", x"48", x"09", x"f0", x"64", x"ab", x"bf", x"5b",
    x"46", x"19", x"f0", x"f5", x"02", x"04", x"26", x"2b",
    x"d7", x"c2", x"00", x"da", x"e4", x"d8", x"d6", x"a9",
    x"05", x"dc", x"f2", x"0e", x"20", x"f9", x"07", x"3d",
    x"31", x"83", x"10", x"00", x"05", x"27", x"25", x"e6",
    x"fb", x"02", x"fc", x"00", x"05", x"fc", x"fd", x"03",
    x"04", x"fc", x"fe", x"fd", x"fd", x"02", x"01", x"ff",
    x"ff", x"03", x"17", x"0c", x"ed", x"4a", x"54", x"41",
    x"10", x"e4", x"f1", x"13", x"ed", x"e2", x"24", x"37",
    x"04", x"fd", x"27", x"3f", x"09", x"19", x"17", x"14",
    x"1f", x"48", x"e9", x"e5", x"f5", x"cc", x"16", x"17",
    x"c7", x"f8", x"1a", x"fb", x"76", x"e4", x"3e", x"37",
    x"25", x"46", x"28", x"1a", x"1d", x"04", x"f3", x"1d",
    x"2b", x"21", x"fd", x"40", x"09", x"f3", x"1c", x"2f",
    x"24", x"02", x"f8", x"f7", x"fd", x"fa", x"0e", x"f9",
    x"14", x"b0", x"de", x"45", x"cd", x"cd", x"19", x"c1",
    x"c7", x"01", x"fd", x"17", x"f5", x"28", x"fc", x"e7",
    x"2e", x"0e", x"17", x"33", x"0c", x"19", x"09", x"e9",
    x"f6", x"6f", x"7e", x"6d", x"f7", x"ef", x"07", x"d9",
    x"27", x"e1", x"d8", x"cb", x"93", x"c3", x"d0", x"e6",
    x"6a", x"de", x"fb", x"32", x"dc", x"ad", x"1d", x"07",
    x"0d", x"1e", x"fe", x"c3", x"8c", x"a5", x"83", x"1f",
    x"72", x"5f", x"c2", x"be", x"08", x"b0", x"d3", x"e5",
    x"02", x"fd", x"fb", x"02", x"fb", x"fd", x"fb", x"fc",
    x"01", x"fb", x"ff", x"f7", x"ff", x"00", x"fa", x"fe",
    x"ff", x"f8", x"fc", x"02", x"03", x"fd", x"fe", x"fa",
    x"02", x"fe", x"06", x"fa", x"fc", x"00", x"f8", x"fb",
    x"fa", x"fb", x"ff", x"fb", x"01", x"00", x"f9", x"00",
    x"fc", x"fe", x"02", x"f7", x"04", x"ff", x"ff", x"fe",
    x"03", x"00", x"ff", x"f7", x"fa", x"fc", x"fe", x"02",
    x"ff", x"03", x"fe", x"f9", x"ff", x"fc", x"00", x"fc",
    x"00", x"00", x"00", x"fd", x"fa", x"fb", x"ff", x"04",
    x"01", x"fe", x"01", x"04", x"01", x"fd", x"fd", x"fe",
    x"fd", x"03", x"fb", x"fb", x"fe", x"f9", x"fe", x"01",
    x"00", x"f7", x"fb", x"02", x"04", x"01", x"ff", x"ff",
    x"04", x"fc", x"04", x"04", x"fe", x"02", x"03", x"02",
    x"04", x"05", x"05", x"ff", x"01", x"05", x"02", x"05",
    x"00", x"fb", x"01", x"fc", x"fc", x"01", x"02", x"fe",
    x"f7", x"fa", x"fd", x"fe", x"fb", x"fb", x"fd", x"fe",
    x"03", x"fd", x"fc", x"fb", x"fe", x"fa", x"fc", x"ff",
    x"fe", x"fd", x"fe", x"01", x"fe", x"01", x"01", x"fd",
    x"fd", x"03", x"fb", x"fa", x"fb", x"01", x"fc", x"ff",
    x"01", x"01", x"ff", x"03", x"03", x"01", x"fb", x"fb",
    x"00", x"04", x"fb", x"fc", x"fc", x"fc", x"04", x"04",
    x"f9", x"fa", x"01", x"fd", x"fe", x"fd", x"fd", x"f9",
    x"01", x"00", x"fd", x"ff", x"ff", x"fd", x"fb", x"ff",
    x"fb", x"fb", x"01", x"00", x"fb", x"fa", x"fc", x"01",
    x"fb", x"00", x"fe", x"f9", x"ff", x"03", x"fd", x"04",
    x"02", x"01", x"fb", x"fe", x"ff", x"03", x"ff", x"fa",
    x"02", x"fa", x"00", x"f9", x"f8", x"01", x"fb", x"fe",
    x"04", x"fc", x"02", x"fd", x"04", x"02", x"02", x"04",
    x"f8", x"00", x"02", x"fe", x"fb", x"fa", x"f6", x"f9",
    x"f9", x"01", x"04", x"fe", x"fd", x"f7", x"f8", x"00",
    x"fd", x"00", x"ff", x"fb", x"02", x"04", x"ff", x"04",
    x"05", x"fc", x"fe", x"00", x"01", x"fb", x"02", x"fd",
    x"fd", x"02", x"fc", x"f9", x"00", x"fb", x"fa", x"fe",
    x"00", x"f8", x"f9", x"01", x"ff", x"01", x"02", x"03",
    x"03", x"ff", x"fa", x"03", x"fb", x"fe", x"01", x"ff",
    x"fd", x"01", x"01", x"fb", x"fd", x"fd", x"fb", x"f8",
    x"ff", x"03", x"fa", x"f7", x"f8", x"01", x"f8", x"f9",
    x"04", x"02", x"03", x"ff", x"fd", x"f9", x"fc", x"f6",
    x"ff", x"fd", x"04", x"fd", x"fc", x"fe", x"00", x"fb",
    x"01", x"03", x"ff", x"f8", x"f9", x"fd", x"fb", x"02",
    x"fd", x"03", x"00", x"f8", x"fb", x"fc", x"fc", x"fb",
    x"00", x"04", x"01", x"ff", x"03", x"03", x"fc", x"00",
    x"fb", x"01", x"03", x"00", x"fb", x"01", x"ff", x"01",
    x"01", x"fd", x"fc", x"ff", x"ff", x"02", x"fb", x"f7",
    x"ff", x"01", x"ff", x"fa", x"fe", x"fc", x"f8", x"fe",
    x"03", x"fe", x"ff", x"04", x"fd", x"03", x"fb", x"fc",
    x"ff", x"fd", x"00", x"fe", x"02", x"f8", x"fa", x"fe",
    x"00", x"fd", x"fb", x"fc", x"03", x"01", x"ff", x"f8",
    x"01", x"fb", x"f9", x"fe", x"03", x"01", x"fc", x"fd",
    x"fb", x"00", x"ff", x"fc", x"fc", x"00", x"03", x"fe",
    x"01", x"00", x"ff", x"f9", x"f7", x"05", x"01", x"fa",
    x"fd", x"fd", x"00", x"fe", x"f7", x"fd", x"03", x"f8",
    x"ff", x"fe", x"fb", x"fb", x"fe", x"fd", x"ff", x"fd",
    x"04", x"fd", x"01", x"01", x"fb", x"fe", x"fc", x"01",
    x"01", x"02", x"00", x"fc", x"fc", x"fb", x"05", x"fe",
    x"00", x"04", x"fa", x"fd", x"fb", x"fe", x"ff", x"02",
    x"03", x"fd", x"ff", x"fa", x"02", x"fb", x"ff", x"fd",
    x"fb", x"fa", x"05", x"ff", x"fb", x"ff", x"fc", x"fb",
    x"f9", x"00", x"fc", x"fa", x"00", x"ff", x"fd", x"01",
    x"04", x"fd", x"fe", x"fc", x"fe", x"02", x"02", x"ff",
    x"01", x"f8", x"fe", x"fa", x"ff", x"fb", x"fe", x"03",
    x"fb", x"03", x"f7", x"00", x"00", x"fe", x"ff", x"fa",
    x"ff", x"00", x"fb", x"fa", x"fd", x"00", x"ff", x"01",
    x"05", x"00", x"03", x"01", x"04", x"fe", x"fe", x"06",
    x"ff", x"fa", x"fc", x"00", x"fc", x"fb", x"01", x"fb",
    x"ff", x"01", x"03", x"ff", x"fe", x"fe", x"f5", x"00",
    x"fb", x"fa", x"f9", x"03", x"02", x"fe", x"fd", x"f7",
    x"f9", x"05", x"f6", x"00", x"fc", x"04", x"03", x"ff",
    x"fa", x"fc", x"f9", x"01", x"01", x"02", x"02", x"f7",
    x"fa", x"f7", x"fd", x"fd", x"fd", x"f6", x"01", x"05",
    x"04", x"01", x"f6", x"fe", x"ff", x"fb", x"00", x"fe",
    x"fd", x"f8", x"fd", x"02", x"fa", x"03", x"04", x"f9",
    x"f5", x"c0", x"be", x"17", x"c6", x"df", x"34", x"44",
    x"27", x"ff", x"04", x"1a", x"46", x"2f", x"18", x"0f",
    x"0b", x"b7", x"ef", x"b1", x"15", x"f2", x"e8", x"d5",
    x"f3", x"d8", x"d4", x"e7", x"e9", x"fd", x"c7", x"d3",
    x"e0", x"d5", x"be", x"cc", x"f5", x"b8", x"d2", x"e6",
    x"02", x"f5", x"fc", x"22", x"07", x"12", x"ee", x"01",
    x"39", x"18", x"c3", x"09", x"14", x"92", x"c7", x"c7",
    x"dd", x"ed", x"da", x"d5", x"12", x"49", x"3f", x"2c",
    x"3b", x"70", x"d1", x"c7", x"b1", x"fa", x"f8", x"0e",
    x"af", x"da", x"d8", x"dc", x"b3", x"8c", x"ef", x"f3",
    x"98", x"0e", x"ee", x"06", x"4f", x"3f", x"34", x"ec",
    x"d5", x"fd", x"cc", x"06", x"19", x"12", x"13", x"1c",
    x"2a", x"20", x"2b", x"bd", x"e8", x"f9", x"ac", x"dc",
    x"05", x"be", x"31", x"31", x"22", x"d8", x"d1", x"06",
    x"d5", x"ba", x"28", x"0b", x"30", x"1f", x"1a", x"45",
    x"ed", x"05", x"42", x"eb", x"00", x"4f", x"41", x"19",
    x"71", x"09", x"fc", x"1b", x"da", x"f6", x"14", x"09",
    x"20", x"0f", x"ff", x"d9", x"fe", x"f0", x"f3", x"05",
    x"2c", x"ef", x"17", x"0b", x"ec", x"05", x"18", x"01",
    x"c9", x"fb", x"fb", x"05", x"fd", x"01", x"03", x"04",
    x"ff", x"04", x"02", x"30", x"29", x"34", x"f8", x"0e",
    x"0c", x"cc", x"c2", x"d7", x"d1", x"e3", x"02", x"e1",
    x"ff", x"d3", x"ce", x"12", x"13", x"17", x"8a", x"0d",
    x"28", x"55", x"e8", x"fb", x"11", x"fb", x"23", x"16",
    x"01", x"27", x"4f", x"f2", x"e7", x"cf", x"2b", x"10",
    x"45", x"1e", x"2f", x"18", x"1b", x"11", x"3b", x"ec",
    x"18", x"d8", x"db", x"28", x"0e", x"14", x"11", x"ff",
    x"df", x"aa", x"d0", x"ef", x"96", x"f4", x"29", x"c0",
    x"d4", x"0c", x"18", x"2e", x"34", x"3b", x"3d", x"48",
    x"1f", x"28", x"fb", x"ee", x"0d", x"10", x"07", x"4d",
    x"f2", x"d7", x"86", x"00", x"fd", x"06", x"07", x"fe",
    x"03", x"ff", x"05", x"fc", x"16", x"d6", x"d3", x"04",
    x"36", x"07", x"da", x"b2", x"c2", x"32", x"de", x"2b",
    x"14", x"28", x"3b", x"4a", x"59", x"49", x"aa", x"06",
    x"cd", x"d9", x"d3", x"e9", x"b6", x"d2", x"c2", x"de",
    x"e9", x"eb", x"d0", x"f8", x"fb", x"12", x"fc", x"3a",
    x"16", x"2e", x"e0", x"1e", x"af", x"fc", x"31", x"08",
    x"ea", x"e4", x"f1", x"0d", x"1b", x"fd", x"03", x"04",
    x"f2", x"22", x"b8", x"2a", x"f0", x"e5", x"ca", x"0c",
    x"17", x"00", x"ee", x"ce", x"d5", x"c0", x"23", x"f4",
    x"18", x"27", x"11", x"06", x"03", x"07", x"05", x"0e",
    x"0a", x"11", x"0a", x"01", x"07", x"d6", x"d0", x"60",
    x"f7", x"09", x"f5", x"3a", x"32", x"0a", x"4a", x"ef",
    x"c7", x"0f", x"e0", x"e7", x"d6", x"db", x"fd", x"a2",
    x"6d", x"89", x"0b", x"f3", x"00", x"0a", x"27", x"36",
    x"00", x"01", x"00", x"00", x"ff", x"03", x"02", x"01",
    x"fe", x"d0", x"b3", x"d4", x"e1", x"eb", x"db", x"d4",
    x"da", x"16", x"f9", x"b5", x"ba", x"d7", x"bc", x"d6",
    x"11", x"09", x"f9", x"d2", x"27", x"18", x"f4", x"fa",
    x"ec", x"05", x"c9", x"ea", x"df", x"c4", x"e1", x"22",
    x"34", x"1d", x"fe", x"24", x"39", x"c1", x"9c", x"1d",
    x"13", x"f4", x"c9", x"fa", x"05", x"02", x"e0", x"c8",
    x"9c", x"30", x"1c", x"08", x"e7", x"fb", x"d1", x"e8",
    x"ee", x"16", x"ea", x"e8", x"f9", x"15", x"0f", x"cb",
    x"fe", x"fb", x"02", x"fa", x"02", x"fd", x"fe", x"fe",
    x"04", x"06", x"03", x"01", x"04", x"06", x"02", x"02",
    x"fa", x"04", x"07", x"e1", x"ed", x"1f", x"41", x"08",
    x"28", x"f0", x"c2", x"ad", x"b9", x"e8", x"fa", x"f8",
    x"1a", x"20", x"e4", x"0d", x"fd", x"f4", x"06", x"21",
    x"38", x"35", x"3f", x"2e", x"20", x"e6", x"28", x"18",
    x"fb", x"f0", x"19", x"e5", x"f9", x"f0", x"01", x"31",
    x"2a", x"1b", x"fd", x"0e", x"2e", x"20", x"11", x"f6",
    x"98", x"a8", x"1f", x"dc", x"f8", x"19", x"55", x"1c",
    x"2d", x"cd", x"cb", x"13", x"d9", x"44", x"18", x"f0",
    x"00", x"eb", x"ff", x"0d", x"23", x"0e", x"de", x"02",
    x"f1", x"12", x"d7", x"eb", x"cd", x"17", x"be", x"d0",
    x"1e", x"39", x"3a", x"32", x"14", x"f6", x"29", x"f5",
    x"07", x"0d", x"bd", x"77", x"ed", x"20", x"e9", x"1c",
    x"b9", x"1a", x"18", x"1b", x"25", x"ae", x"c1", x"b7",
    x"1e", x"f4", x"0f", x"16", x"1f", x"0e", x"03", x"b6",
    x"c2", x"fa", x"9d", x"7b", x"18", x"c1", x"b4", x"ad",
    x"02", x"09", x"f3", x"dc", x"b4", x"02", x"05", x"fe",
    x"13", x"04", x"f6", x"2c", x"2d", x"f4", x"30", x"4e",
    x"d3", x"b8", x"f5", x"1c", x"fd", x"ec", x"19", x"18",
    x"fe", x"02", x"e2", x"e8", x"d9", x"07", x"eb", x"d2",
    x"fe", x"f2", x"d9", x"11", x"1d", x"01", x"cb", x"ba",
    x"e4", x"e1", x"1b", x"ed", x"e4", x"17", x"0f", x"38",
    x"42", x"04", x"5a", x"2e", x"fb", x"d0", x"ea", x"13",
    x"fa", x"f4", x"e7", x"ce", x"f4", x"e7", x"cf", x"1d",
    x"d8", x"e5", x"ec", x"ae", x"0e", x"b7", x"8d", x"0f",
    x"f0", x"12", x"e4", x"dc", x"bb", x"ee", x"ec", x"bb",
    x"2a", x"13", x"05", x"1f", x"01", x"f5", x"f6", x"e7",
    x"e1", x"31", x"47", x"4c", x"d4", x"b1", x"fa", x"e0",
    x"d9", x"f6", x"10", x"ee", x"fd", x"fe", x"2a", x"39",
    x"4f", x"0f", x"f5", x"e3", x"cd", x"f0", x"bb", x"d0",
    x"f4", x"f5", x"f5", x"fb", x"28", x"30", x"1f", x"14",
    x"4c", x"22", x"3f", x"12", x"d2", x"e3", x"cc", x"7f",
    x"e5", x"e1", x"d7", x"04", x"fc", x"b2", x"3a", x"10",
    x"12", x"0a", x"c2", x"da", x"e3", x"d6", x"da", x"34",
    x"1b", x"e5", x"33", x"24", x"35", x"21", x"1e", x"28",
    x"2d", x"1b", x"78", x"2c", x"2e", x"47", x"27", x"eb",
    x"db", x"fa", x"ff", x"ff", x"01", x"00", x"fc", x"01",
    x"fc", x"04", x"cd", x"d5", x"06", x"6d", x"1e", x"b9",
    x"d2", x"e4", x"ef", x"de", x"e9", x"0e", x"c8", x"c2",
    x"03", x"cb", x"e8", x"bc", x"e3", x"ee", x"05", x"fb",
    x"f0", x"0f", x"f9", x"16", x"d2", x"e0", x"f7", x"16",
    x"e3", x"de", x"dd", x"d9", x"6c", x"61", x"f1", x"00",
    x"16", x"2c", x"23", x"21", x"36", x"fb", x"b8", x"f9",
    x"20", x"0d", x"0f", x"1c", x"17", x"50", x"30", x"22",
    x"c9", x"bd", x"cb", x"08", x"05", x"f6", x"fa", x"2d",
    x"03", x"e8", x"f2", x"0d", x"0e", x"38", x"3a", x"64",
    x"59", x"2c", x"e5", x"fb", x"15", x"e7", x"fd", x"05",
    x"e0", x"7c", x"a2", x"fe", x"fa", x"f3", x"fb", x"fa",
    x"ff", x"fc", x"07", x"fc", x"1c", x"4c", x"3e", x"17",
    x"29", x"26", x"ff", x"17", x"2d", x"fe", x"25", x"63",
    x"f9", x"0b", x"3f", x"1c", x"27", x"20", x"ec", x"e9",
    x"ed", x"e7", x"e1", x"f9", x"a1", x"bd", x"c2", x"0e",
    x"01", x"1b", x"12", x"e4", x"05", x"fe", x"d3", x"ec",
    x"2f", x"44", x"e7", x"13", x"26", x"39", x"21", x"2e",
    x"1b", x"fe", x"e1", x"35", x"ed", x"05", x"17", x"16",
    x"0d", x"3b", x"df", x"ea", x"b2", x"e5", x"e8", x"ea",
    x"f9", x"f1", x"cf", x"14", x"1c", x"fa", x"ec", x"01",
    x"08", x"d0", x"1d", x"1a", x"13", x"fd", x"02", x"0f",
    x"03", x"f9", x"14", x"02", x"f8", x"03", x"06", x"1b",
    x"25", x"0e", x"22", x"00", x"10", x"fe", x"29", x"09",
    x"3c", x"3e", x"f5", x"05", x"73", x"fb", x"ef", x"22",
    x"fe", x"fd", x"1d", x"01", x"d0", x"01", x"d1", x"a5",
    x"fd", x"01", x"05", x"02", x"fe", x"05", x"fe", x"ff",
    x"06", x"d4", x"ff", x"fc", x"00", x"e4", x"f8", x"f4",
    x"e2", x"e2", x"01", x"f2", x"0c", x"f8", x"ee", x"04",
    x"d7", x"e7", x"ec", x"c5", x"ec", x"fc", x"04", x"f2",
    x"0b", x"f4", x"1f", x"2e", x"fb", x"ef", x"c2", x"d9",
    x"f2", x"24", x"c3", x"0c", x"0d", x"27", x"0b", x"3c",
    x"0d", x"0d", x"fe", x"2a", x"23", x"13", x"cc", x"f1",
    x"1c", x"b3", x"c8", x"0e", x"ee", x"f3", x"13", x"c3",
    x"b0", x"e2", x"fb", x"d1", x"ef", x"ed", x"e3", x"b0",
    x"01", x"01", x"04", x"f5", x"fd", x"ff", x"04", x"02",
    x"06", x"01", x"00", x"fc", x"01", x"06", x"fc", x"00",
    x"fa", x"02", x"f1", x"32", x"3a", x"29", x"31", x"2d",
    x"59", x"39", x"60", x"2f", x"fe", x"fd", x"01", x"06",
    x"da", x"16", x"b8", x"85", x"b9", x"b3", x"21", x"cb",
    x"f3", x"41", x"aa", x"ce", x"22", x"15", x"1e", x"0c",
    x"df", x"e2", x"f7", x"06", x"d9", x"04", x"21", x"fb",
    x"f0", x"68", x"c1", x"05", x"ba", x"da", x"01", x"c1",
    x"d2", x"e6", x"32", x"fa", x"07", x"f8", x"bb", x"af",
    x"00", x"17", x"01", x"0b", x"fa", x"0a", x"37", x"28",
    x"1c", x"d6", x"fb", x"22", x"ff", x"2b", x"49", x"ef",
    x"11", x"33", x"36", x"2b", x"b9", x"38", x"22", x"15",
    x"46", x"4b", x"46", x"e9", x"f4", x"19", x"e3", x"db",
    x"cd", x"fa", x"c3", x"ca", x"3b", x"2f", x"14", x"cf",
    x"18", x"14", x"36", x"23", x"09", x"fa", x"23", x"11",
    x"27", x"0b", x"24", x"ed", x"29", x"0f", x"45", x"2b",
    x"0e", x"1d", x"0e", x"fb", x"18", x"f6", x"1c", x"d4",
    x"d4", x"14", x"e8", x"f5", x"ff", x"40", x"09", x"09",
    x"fc", x"00", x"04", x"fa", x"03", x"fe", x"fa", x"00",
    x"05", x"fb", x"fe", x"00", x"fa", x"fc", x"f8", x"fa",
    x"00", x"fe", x"fa", x"03", x"02", x"fd", x"fa", x"ff",
    x"f8", x"fa", x"00", x"fa", x"fb", x"00", x"00", x"fb",
    x"00", x"fd", x"ff", x"ff", x"02", x"00", x"fa", x"00",
    x"ff", x"02", x"fc", x"03", x"00", x"fc", x"fe", x"fc",
    x"00", x"00", x"f9", x"f7", x"fd", x"fa", x"fe", x"fe",
    x"fb", x"fc", x"03", x"fd", x"02", x"fc", x"fc", x"00",
    x"04", x"03", x"02", x"fb", x"03", x"fb", x"ff", x"ff",
    x"03", x"fa", x"fd", x"fe", x"fe", x"fb", x"fa", x"fe",
    x"02", x"fb", x"01", x"02", x"ff", x"fa", x"fc", x"fc",
    x"fb", x"fa", x"04", x"fd", x"fb", x"03", x"fc", x"03",
    x"fe", x"fa", x"01", x"02", x"fd", x"03", x"03", x"05",
    x"05", x"ff", x"fa", x"ff", x"00", x"fe", x"fb", x"fd",
    x"fb", x"01", x"04", x"ff", x"fa", x"ff", x"fb", x"ff",
    x"fb", x"02", x"02", x"f7", x"fc", x"fe", x"fe", x"fb",
    x"05", x"02", x"fe", x"fc", x"ff", x"01", x"01", x"04",
    x"ff", x"fb", x"04", x"fb", x"fe", x"02", x"fb", x"01",
    x"00", x"00", x"03", x"fb", x"fe", x"fa", x"ff", x"ff",
    x"ff", x"fc", x"ff", x"03", x"01", x"05", x"fe", x"00",
    x"fd", x"03", x"04", x"04", x"01", x"fa", x"01", x"01",
    x"fc", x"fb", x"00", x"fe", x"ff", x"fe", x"f9", x"fb",
    x"f8", x"fa", x"00", x"04", x"fd", x"ff", x"fe", x"fe",
    x"f8", x"ff", x"f9", x"f8", x"01", x"fa", x"05", x"ff",
    x"02", x"ff", x"fd", x"03", x"fe", x"fd", x"03", x"ff",
    x"00", x"02", x"02", x"01", x"01", x"fe", x"04", x"01",
    x"fb", x"fe", x"fc", x"fe", x"fb", x"fa", x"fe", x"fd",
    x"ff", x"01", x"fe", x"03", x"00", x"04", x"fc", x"fc",
    x"f7", x"01", x"f7", x"02", x"00", x"00", x"ff", x"fc",
    x"00", x"fd", x"00", x"03", x"fa", x"f9", x"f8", x"ff",
    x"fa", x"fb", x"fa", x"02", x"02", x"fe", x"fb", x"04",
    x"04", x"04", x"ff", x"04", x"01", x"fb", x"04", x"02",
    x"fc", x"04", x"fe", x"f9", x"01", x"fc", x"fd", x"f9",
    x"fd", x"fe", x"fd", x"02", x"fc", x"fa", x"00", x"01",
    x"ff", x"fe", x"01", x"01", x"03", x"fc", x"01", x"04",
    x"03", x"02", x"fd", x"01", x"f8", x"fa", x"00", x"fd",
    x"fe", x"04", x"fb", x"fa", x"01", x"fb", x"03", x"ff",
    x"fe", x"01", x"fa", x"f9", x"00", x"ff", x"f9", x"fe",
    x"fc", x"fb", x"ff", x"00", x"fd", x"01", x"fd", x"00",
    x"fb", x"02", x"fd", x"fa", x"02", x"fe", x"f9", x"02",
    x"fe", x"02", x"04", x"04", x"fd", x"01", x"00", x"fb",
    x"00", x"ff", x"fe", x"ff", x"fb", x"02", x"fd", x"04",
    x"fb", x"fe", x"fd", x"fc", x"fc", x"f9", x"03", x"fc",
    x"fc", x"04", x"ff", x"fb", x"04", x"ff", x"ff", x"02",
    x"fc", x"fe", x"f9", x"fc", x"fd", x"04", x"fc", x"01",
    x"05", x"fc", x"04", x"fc", x"fe", x"05", x"04", x"01",
    x"05", x"fc", x"03", x"02", x"fc", x"ff", x"00", x"fe",
    x"fb", x"ff", x"02", x"fc", x"fc", x"fe", x"fd", x"fd",
    x"fb", x"ff", x"fd", x"ff", x"ff", x"03", x"fb", x"fb",
    x"f8", x"03", x"fe", x"f9", x"fd", x"03", x"fc", x"fb",
    x"00", x"fb", x"00", x"fc", x"fa", x"fc", x"03", x"fa",
    x"ff", x"03", x"00", x"f9", x"fe", x"fc", x"01", x"00",
    x"ff", x"fc", x"00", x"fc", x"fc", x"fa", x"02", x"01",
    x"fc", x"00", x"fd", x"fb", x"fa", x"fb", x"01", x"f9",
    x"01", x"02", x"fc", x"fe", x"02", x"fe", x"02", x"04",
    x"fc", x"ff", x"04", x"00", x"fe", x"fe", x"03", x"05",
    x"fc", x"02", x"fc", x"fe", x"01", x"fb", x"fb", x"ff",
    x"fc", x"ff", x"f9", x"02", x"f9", x"fc", x"f9", x"fb",
    x"fc", x"f8", x"01", x"00", x"fb", x"fe", x"fe", x"03",
    x"f7", x"fb", x"01", x"fa", x"f7", x"fc", x"01", x"fd",
    x"f7", x"ff", x"f9", x"00", x"fa", x"03", x"fd", x"01",
    x"fe", x"02", x"04", x"fb", x"fb", x"fc", x"01", x"00",
    x"03", x"fc", x"ff", x"fe", x"fe", x"04", x"03", x"01",
    x"02", x"01", x"fb", x"04", x"fc", x"03", x"fc", x"03",
    x"01", x"fc", x"fd", x"01", x"fe", x"fe", x"fc", x"fe",
    x"02", x"fd", x"fd", x"03", x"05", x"fd", x"02", x"fb",
    x"03", x"fb", x"f8", x"03", x"ff", x"01", x"f8", x"01",
    x"fc", x"f7", x"f7", x"00", x"04", x"04", x"ff", x"02",
    x"fa", x"03", x"f9", x"fd", x"01", x"02", x"01", x"01",
    x"fe", x"f8", x"fa", x"fd", x"f8", x"00", x"00", x"02",
    x"fd", x"ff", x"01", x"01", x"f9", x"fe", x"fa", x"fe",
    x"01", x"00", x"fb", x"ff", x"02", x"00", x"00", x"02",
    x"d4", x"bc", x"b3", x"28", x"fe", x"04", x"1d", x"24",
    x"25", x"fe", x"f6", x"d4", x"e7", x"10", x"19", x"c4",
    x"03", x"19", x"c9", x"b6", x"61", x"ae", x"9a", x"a0",
    x"d6", x"a0", x"b0", x"31", x"1b", x"2a", x"15", x"ee",
    x"f8", x"e2", x"c4", x"ed", x"b1", x"be", x"d2", x"ba",
    x"cb", x"b9", x"aa", x"b6", x"b7", x"d0", x"36", x"03",
    x"c2", x"04", x"24", x"d9", x"d3", x"ea", x"f9", x"06",
    x"fa", x"03", x"05", x"19", x"0c", x"c7", x"d1", x"14",
    x"18", x"fc", x"1b", x"04", x"22", x"fb", x"06", x"11",
    x"ac", x"03", x"b4", x"dc", x"c4", x"f9", x"dd", x"e1",
    x"ff", x"bd", x"17", x"28", x"19", x"30", x"15", x"2e",
    x"39", x"21", x"19", x"c0", x"78", x"d5", x"83", x"9e",
    x"61", x"05", x"e2", x"4b", x"db", x"12", x"f8", x"f2",
    x"04", x"2a", x"fe", x"00", x"0f", x"b3", x"d6", x"14",
    x"e1", x"b5", x"ed", x"06", x"f5", x"b4", x"d0", x"b4",
    x"df", x"08", x"c0", x"0f", x"06", x"7f", x"12", x"d0",
    x"ad", x"12", x"1c", x"e1", x"02", x"f3", x"00", x"ac",
    x"a5", x"14", x"b2", x"ce", x"f7", x"e4", x"af", x"09",
    x"15", x"1c", x"f5", x"e5", x"0f", x"12", x"f1", x"08",
    x"39", x"05", x"ff", x"fd", x"ff", x"fe", x"00", x"ff",
    x"ff", x"fe", x"a3", x"a1", x"01", x"24", x"cf", x"4a",
    x"07", x"1a", x"35", x"f4", x"ea", x"1b", x"eb", x"10",
    x"1f", x"43", x"26", x"15", x"12", x"e3", x"9d", x"ea",
    x"ec", x"7b", x"ea", x"e3", x"08", x"d2", x"cf", x"a2",
    x"c4", x"f9", x"e1", x"11", x"1d", x"0a", x"12", x"23",
    x"dd", x"1c", x"2d", x"33", x"c8", x"13", x"31", x"da",
    x"e7", x"e3", x"09", x"e8", x"fc", x"f0", x"02", x"4c",
    x"5a", x"eb", x"bd", x"f8", x"30", x"25", x"e9", x"22",
    x"2b", x"f5", x"a3", x"6e", x"e4", x"ce", x"a9", x"16",
    x"52", x"4c", x"ae", x"d5", x"d8", x"98", x"de", x"e6",
    x"33", x"25", x"1f", x"0c", x"06", x"05", x"fa", x"0a",
    x"fb", x"01", x"08", x"04", x"cf", x"ec", x"f4", x"b0",
    x"b7", x"bc", x"fd", x"1b", x"1b", x"09", x"ef", x"fe",
    x"f2", x"cc", x"b9", x"d6", x"bd", x"c7", x"df", x"13",
    x"f7", x"40", x"2c", x"94", x"11", x"27", x"34", x"07",
    x"d1", x"20", x"d5", x"f6", x"0b", x"fa", x"fc", x"f9",
    x"d1", x"8e", x"a7", x"01", x"e9", x"7c", x"0b", x"fd",
    x"ef", x"1e", x"c8", x"da", x"f8", x"00", x"f7", x"1d",
    x"19", x"d6", x"66", x"b2", x"e4", x"1a", x"f1", x"07",
    x"26", x"00", x"19", x"c8", x"00", x"fd", x"45", x"1c",
    x"e8", x"41", x"29", x"24", x"fd", x"08", x"01", x"03",
    x"0d", x"04", x"01", x"00", x"09", x"1a", x"a1", x"6d",
    x"37", x"d5", x"92", x"d0", x"df", x"b4", x"74", x"ce",
    x"ae", x"fc", x"d4", x"f4", x"06", x"e6", x"db", x"48",
    x"24", x"12", x"01", x"eb", x"ea", x"ef", x"a1", x"88",
    x"04", x"fd", x"fd", x"03", x"01", x"fe", x"02", x"01",
    x"00", x"25", x"ce", x"c9", x"17", x"97", x"78", x"2c",
    x"12", x"03", x"22", x"f7", x"1b", x"1e", x"f8", x"c0",
    x"eb", x"23", x"07", x"12", x"c8", x"d1", x"2c", x"23",
    x"c7", x"4f", x"18", x"32", x"1b", x"22", x"e2", x"f3",
    x"b7", x"21", x"24", x"04", x"cd", x"ea", x"df", x"fc",
    x"10", x"e9", x"ee", x"f2", x"0e", x"23", x"d0", x"09",
    x"fd", x"0a", x"0b", x"1b", x"33", x"14", x"27", x"df",
    x"15", x"dc", x"dc", x"2c", x"32", x"2b", x"16", x"17",
    x"03", x"04", x"03", x"fd", x"fc", x"01", x"03", x"01",
    x"00", x"03", x"03", x"00", x"05", x"ff", x"02", x"03",
    x"fc", x"05", x"f8", x"f7", x"e4", x"1c", x"2f", x"10",
    x"dd", x"e8", x"f8", x"01", x"d8", x"8d", x"2d", x"3f",
    x"89", x"12", x"26", x"e2", x"d3", x"d5", x"06", x"c1",
    x"ea", x"42", x"f1", x"fe", x"0a", x"ef", x"1e", x"0c",
    x"31", x"28", x"18", x"eb", x"11", x"10", x"30", x"fe",
    x"ea", x"b8", x"de", x"fd", x"d9", x"aa", x"21", x"37",
    x"f9", x"e4", x"1b", x"f5", x"f4", x"02", x"c8", x"d2",
    x"17", x"13", x"dd", x"30", x"df", x"f2", x"32", x"c7",
    x"d2", x"23", x"26", x"2d", x"12", x"21", x"42", x"e0",
    x"e7", x"2d", x"11", x"0e", x"f2", x"1d", x"0c", x"1f",
    x"09", x"d9", x"e0", x"1d", x"0e", x"04", x"25", x"eb",
    x"d7", x"04", x"1b", x"1e", x"fb", x"43", x"fb", x"07",
    x"65", x"18", x"15", x"3d", x"3a", x"ea", x"13", x"28",
    x"07", x"e9", x"24", x"0c", x"f8", x"d5", x"3b", x"22",
    x"fd", x"fc", x"0b", x"0f", x"e0", x"ee", x"23", x"31",
    x"d1", x"98", x"24", x"12", x"52", x"00", x"07", x"42",
    x"43", x"1f", x"40", x"46", x"08", x"d2", x"ec", x"fb",
    x"44", x"c9", x"11", x"24", x"00", x"23", x"fd", x"cd",
    x"ad", x"91", x"ea", x"aa", x"ba", x"b2", x"ac", x"c8",
    x"df", x"0d", x"02", x"e9", x"d7", x"fb", x"de", x"e3",
    x"10", x"25", x"0c", x"0f", x"d0", x"cb", x"e9", x"c6",
    x"ce", x"f4", x"b5", x"cb", x"f1", x"ad", x"f1", x"08",
    x"bb", x"f2", x"02", x"d9", x"fe", x"e8", x"eb", x"1a",
    x"fa", x"f8", x"e3", x"d8", x"d8", x"fe", x"68", x"c7",
    x"0a", x"05", x"11", x"1f", x"2a", x"27", x"1f", x"f6",
    x"bc", x"ea", x"fc", x"20", x"22", x"19", x"2c", x"2c",
    x"ef", x"ea", x"ef", x"13", x"08", x"1f", x"f6", x"f0",
    x"0b", x"e7", x"f4", x"de", x"ce", x"44", x"e9", x"f1",
    x"3b", x"f4", x"2b", x"3b", x"e7", x"c1", x"2c", x"ca",
    x"c1", x"ab", x"1e", x"36", x"0f", x"11", x"fa", x"ff",
    x"df", x"c3", x"c0", x"a8", x"a1", x"b6", x"fa", x"fb",
    x"12", x"f5", x"ef", x"f4", x"03", x"43", x"ee", x"cf",
    x"e1", x"e7", x"da", x"fb", x"fd", x"03", x"02", x"a8",
    x"ba", x"a7", x"86", x"75", x"be", x"91", x"b7", x"27",
    x"f1", x"13", x"29", x"14", x"09", x"32", x"ea", x"d7",
    x"fa", x"03", x"ff", x"04", x"fd", x"fd", x"fc", x"ff",
    x"00", x"05", x"bf", x"b6", x"c6", x"f4", x"33", x"f5",
    x"2b", x"00", x"11", x"ec", x"12", x"18", x"0d", x"22",
    x"56", x"0c", x"3d", x"20", x"d9", x"de", x"bd", x"df",
    x"ec", x"15", x"05", x"f0", x"17", x"ce", x"0f", x"f6",
    x"1a", x"37", x"2a", x"17", x"29", x"0d", x"0b", x"1c",
    x"2e", x"e4", x"21", x"03", x"c2", x"cc", x"45", x"ab",
    x"e1", x"13", x"fa", x"17", x"31", x"dd", x"f5", x"02",
    x"5d", x"12", x"01", x"b7", x"06", x"e9", x"fb", x"c7",
    x"e2", x"d4", x"be", x"fb", x"0d", x"f8", x"26", x"ed",
    x"e7", x"f5", x"d7", x"fa", x"13", x"3c", x"41", x"3b",
    x"fd", x"51", x"15", x"04", x"00", x"f9", x"06", x"fd",
    x"02", x"fd", x"fe", x"fb", x"99", x"cc", x"e5", x"12",
    x"06", x"10", x"30", x"08", x"08", x"0e", x"10", x"17",
    x"f8", x"0a", x"07", x"22", x"37", x"06", x"e6", x"b7",
    x"a3", x"0f", x"02", x"05", x"f0", x"0a", x"0d", x"d3",
    x"e5", x"ea", x"f6", x"fc", x"15", x"ea", x"08", x"fc",
    x"02", x"0d", x"dc", x"15", x"0a", x"d0", x"02", x"e9",
    x"f7", x"b9", x"ff", x"23", x"3c", x"32", x"24", x"1d",
    x"f5", x"fd", x"19", x"0b", x"d1", x"20", x"eb", x"94",
    x"05", x"cb", x"74", x"32", x"20", x"f7", x"33", x"37",
    x"06", x"7e", x"3c", x"14", x"f7", x"02", x"07", x"01",
    x"07", x"03", x"01", x"ff", x"07", x"41", x"cd", x"90",
    x"01", x"fe", x"27", x"20", x"2a", x"2e", x"66", x"c3",
    x"83", x"51", x"ce", x"d8", x"b1", x"05", x"0d", x"34",
    x"d4", x"92", x"e0", x"ca", x"f9", x"a0", x"f1", x"02",
    x"04", x"fd", x"fb", x"fe", x"00", x"01", x"05", x"01",
    x"fc", x"c1", x"cd", x"91", x"c5", x"dd", x"ee", x"3e",
    x"23", x"31", x"d1", x"a9", x"dc", x"31", x"28", x"31",
    x"62", x"43", x"4d", x"09", x"d3", x"de", x"36", x"3e",
    x"18", x"3f", x"1b", x"ed", x"cf", x"25", x"f1", x"d9",
    x"ea", x"22", x"d8", x"e5", x"00", x"14", x"ed", x"1b",
    x"1b", x"13", x"fa", x"19", x"1d", x"fc", x"de", x"29",
    x"03", x"10", x"eb", x"cd", x"f1", x"04", x"f6", x"17",
    x"3c", x"14", x"1a", x"03", x"04", x"2d", x"f5", x"c4",
    x"02", x"01", x"01", x"00", x"fc", x"fc", x"04", x"fc",
    x"fc", x"06", x"ff", x"fc", x"fa", x"fc", x"fc", x"03",
    x"06", x"01", x"39", x"16", x"2b", x"ee", x"1f", x"2d",
    x"d9", x"b5", x"ab", x"23", x"73", x"a1", x"23", x"f4",
    x"df", x"35", x"04", x"06", x"f1", x"e3", x"2b", x"de",
    x"b9", x"de", x"f5", x"05", x"1e", x"f4", x"f3", x"f3",
    x"0e", x"09", x"fb", x"d4", x"d6", x"c1", x"2b", x"1a",
    x"df", x"3b", x"10", x"da", x"22", x"26", x"14", x"5b",
    x"f2", x"19", x"fe", x"c7", x"c7", x"bc", x"0e", x"01",
    x"0f", x"08", x"b9", x"2a", x"f4", x"cf", x"fb", x"1b",
    x"e8", x"d4", x"06", x"f3", x"1f", x"f0", x"1a", x"bb",
    x"99", x"cf", x"de", x"24", x"e7", x"c8", x"c7", x"90",
    x"d4", x"08", x"1e", x"f8", x"ff", x"04", x"d7", x"e6",
    x"f6", x"e0", x"f6", x"a7", x"1b", x"1b", x"02", x"3c",
    x"49", x"16", x"22", x"2a", x"15", x"0c", x"14", x"34",
    x"35", x"47", x"2f", x"18", x"0c", x"ef", x"0a", x"f3",
    x"0e", x"1c", x"0d", x"0b", x"f5", x"e2", x"9f", x"14",
    x"1e", x"4d", x"d5", x"07", x"e4", x"ed", x"c7", x"db",
    x"28", x"10", x"9e", x"09", x"20", x"cb", x"08", x"0a",
    x"f0", x"04", x"e2", x"34", x"a2", x"d4", x"fb", x"26",
    x"22", x"27", x"ea", x"dc", x"b5", x"8b", x"d0", x"a2",
    x"8e", x"ba", x"e9", x"fd", x"ea", x"0e", x"08", x"23",
    x"49", x"11", x"0e", x"0c", x"e7", x"0e", x"05", x"dc",
    x"ce", x"c8", x"b1", x"c2", x"02", x"f9", x"32", x"25",
    x"f1", x"01", x"00", x"3e", x"19", x"fe", x"f0", x"15",
    x"fd", x"25", x"43", x"f6", x"fe", x"2b", x"2c", x"ea",
    x"94", x"ec", x"33", x"f4", x"16", x"e9", x"ed", x"29",
    x"12", x"e3", x"db", x"18", x"fe", x"30", x"bc", x"df",
    x"f3", x"d9", x"c7", x"cd", x"98", x"c2", x"1b", x"ba",
    x"90", x"20", x"2c", x"de", x"3e", x"2c", x"c4", x"0b",
    x"f7", x"f6", x"0a", x"e6", x"1e", x"f6", x"49", x"19",
    x"00", x"19", x"1c", x"fc", x"e4", x"05", x"02", x"56",
    x"fa", x"f1", x"fc", x"ed", x"ee", x"bd", x"c7", x"19",
    x"ee", x"f3", x"1e", x"f4", x"e5", x"ce", x"0f", x"0d",
    x"2d", x"72", x"be", x"e7", x"d4", x"e3", x"de", x"c4",
    x"e3", x"dd", x"f1", x"f9", x"e4", x"39", x"23", x"0c",
    x"1e", x"02", x"07", x"f5", x"2b", x"2d", x"c6", x"b9",
    x"22", x"02", x"ff", x"03", x"06", x"fd", x"fb", x"01",
    x"fe", x"fd", x"fa", x"f1", x"46", x"b2", x"90", x"e1",
    x"01", x"14", x"08", x"b3", x"0e", x"0b", x"bc", x"fe",
    x"35", x"03", x"1a", x"16", x"0d", x"0b", x"25", x"35",
    x"0a", x"e1", x"3d", x"41", x"e7", x"fa", x"08", x"15",
    x"bb", x"f9", x"24", x"d0", x"c7", x"d9", x"21", x"0c",
    x"28", x"d1", x"f3", x"e2", x"ff", x"b7", x"c2", x"d4",
    x"e9", x"1c", x"b0", x"ea", x"ea", x"23", x"c4", x"d4",
    x"14", x"32", x"06", x"40", x"0c", x"c0", x"bb", x"13",
    x"b7", x"db", x"e1", x"42", x"1e", x"17", x"20", x"2e",
    x"40", x"12", x"d9", x"15", x"0a", x"b1", x"00", x"20",
    x"1b", x"45", x"0d", x"01", x"02", x"fa", x"00", x"05",
    x"fc", x"02", x"01", x"03", x"30", x"10", x"09", x"fd",
    x"e7", x"05", x"ff", x"1b", x"ee", x"f9", x"30", x"37",
    x"e7", x"1f", x"1a", x"08", x"15", x"06", x"c4", x"d6",
    x"fc", x"00", x"be", x"9f", x"c6", x"92", x"c5", x"28",
    x"d5", x"f2", x"f0", x"e7", x"f5", x"d4", x"eb", x"41",
    x"09", x"25", x"e7", x"2f", x"2b", x"d0", x"17", x"2b",
    x"78", x"9e", x"e0", x"07", x"da", x"86", x"fd", x"1f",
    x"0b", x"3a", x"24", x"47", x"2f", x"f8", x"34", x"07",
    x"e0", x"15", x"e2", x"0e", x"2f", x"ee", x"2d", x"bd",
    x"22", x"da", x"fd", x"02", x"08", x"01", x"00", x"06",
    x"fd", x"ff", x"03", x"01", x"fd", x"07", x"2a", x"17",
    x"00", x"26", x"35", x"e1", x"e5", x"fb", x"3e", x"c2",
    x"c3", x"7d", x"d2", x"ab", x"43", x"ec", x"ad", x"13",
    x"25", x"cd", x"42", x"0a", x"b5", x"29", x"09", x"d2",
    x"fb", x"00", x"04", x"fc", x"fe", x"00", x"fc", x"fc",
    x"04", x"ed", x"b7", x"b4", x"bb", x"e5", x"ea", x"dc",
    x"c7", x"e6", x"e0", x"20", x"e5", x"90", x"1d", x"3c",
    x"f4", x"e1", x"2b", x"1d", x"d4", x"e8", x"03", x"74",
    x"c8", x"07", x"49", x"9b", x"d9", x"c1", x"fe", x"04",
    x"f4", x"1b", x"f3", x"c6", x"f0", x"37", x"15", x"39",
    x"00", x"de", x"e6", x"d6", x"f4", x"b1", x"f4", x"59",
    x"24", x"c3", x"07", x"12", x"e5", x"d6", x"fd", x"16",
    x"11", x"21", x"f7", x"10", x"06", x"bf", x"f1", x"d0",
    x"00", x"fe", x"03", x"fe", x"ff", x"fd", x"02", x"ff",
    x"05", x"fd", x"fa", x"01", x"fe", x"fb", x"01", x"01",
    x"fd", x"04", x"79", x"26", x"34", x"ee", x"0f", x"38",
    x"c3", x"ff", x"eb", x"31", x"41", x"13", x"14", x"03",
    x"9b", x"ff", x"f6", x"a7", x"dc", x"db", x"16", x"9b",
    x"d4", x"ba", x"00", x"c5", x"01", x"d2", x"ec", x"f5",
    x"e8", x"02", x"36", x"ea", x"f9", x"3c", x"1c", x"13",
    x"f6", x"0d", x"0f", x"f9", x"18", x"01", x"d5", x"10",
    x"21", x"20", x"33", x"12", x"08", x"ef", x"17", x"f7",
    x"1b", x"3c", x"f2", x"01", x"29", x"e6", x"2e", x"01",
    x"e5", x"f7", x"20", x"2a", x"e0", x"15", x"46", x"c4",
    x"44", x"47", x"d8", x"07", x"d4", x"ff", x"05", x"16",
    x"07", x"11", x"2c", x"ec", x"20", x"17", x"f5", x"01",
    x"c4", x"0b", x"ec", x"b8", x"e3", x"e1", x"00", x"e7",
    x"38", x"32", x"d3", x"ed", x"f2", x"1f", x"17", x"13",
    x"f5", x"ed", x"f8", x"e2", x"e7", x"29", x"f4", x"ff",
    x"f2", x"3e", x"02", x"11", x"34", x"fa", x"ed", x"ff",
    x"34", x"1c", x"08", x"fc", x"e6", x"f1", x"0b", x"15",
    x"e6", x"cc", x"9b", x"05", x"ba", x"c2", x"0f", x"f8",
    x"04", x"0e", x"e9", x"d0", x"ac", x"1a", x"05", x"ec",
    x"03", x"11", x"f1", x"f0", x"d2", x"fd", x"0d", x"14",
    x"dc", x"f0", x"dc", x"dd", x"d9", x"ed", x"15", x"b3",
    x"de", x"3d", x"25", x"cc", x"f7", x"e3", x"df", x"1c",
    x"11", x"54", x"55", x"57", x"46", x"34", x"17", x"07",
    x"10", x"ff", x"e4", x"bf", x"eb", x"c1", x"0b", x"f9",
    x"f5", x"cc", x"e9", x"eb", x"f9", x"21", x"15", x"2e",
    x"21", x"1f", x"eb", x"ee", x"f5", x"c2", x"d4", x"e0",
    x"14", x"08", x"f8", x"15", x"18", x"04", x"0f", x"06",
    x"1c", x"1f", x"3e", x"3f", x"ed", x"f8", x"fb", x"05",
    x"e9", x"dd", x"b7", x"b6", x"d9", x"42", x"bb", x"d6",
    x"12", x"d4", x"e5", x"f5", x"13", x"44", x"2a", x"e1",
    x"f4", x"eb", x"af", x"b3", x"d2", x"25", x"fa", x"e7",
    x"e2", x"e1", x"00", x"ea", x"e6", x"db", x"97", x"96",
    x"46", x"21", x"bf", x"19", x"19", x"34", x"1e", x"4c",
    x"34", x"21", x"3f", x"40", x"65", x"39", x"3f", x"f9",
    x"1a", x"3a", x"ec", x"f7", x"1a", x"20", x"fe", x"cd",
    x"e2", x"06", x"11", x"da", x"f4", x"17", x"9d", x"d0",
    x"e4", x"fc", x"02", x"03", x"ff", x"03", x"00", x"fe",
    x"01", x"fe", x"0e", x"eb", x"dd", x"26", x"20", x"ec",
    x"ed", x"d7", x"d7", x"19", x"06", x"c8", x"fa", x"0b",
    x"db", x"0c", x"1c", x"1c", x"06", x"e4", x"f8", x"ef",
    x"f4", x"ff", x"a8", x"ee", x"21", x"dc", x"0e", x"05",
    x"e8", x"ef", x"e8", x"d8", x"fe", x"15", x"01", x"ff",
    x"f1", x"f1", x"df", x"b1", x"bc", x"ec", x"23", x"f9",
    x"0b", x"e7", x"fb", x"04", x"fc", x"18", x"12", x"f1",
    x"ef", x"af", x"d3", x"0f", x"16", x"23", x"82", x"20",
    x"1b", x"28", x"1e", x"d4", x"f2", x"1b", x"e7", x"cd",
    x"24", x"fd", x"20", x"ef", x"f1", x"27", x"0d", x"ec",
    x"a2", x"ed", x"e5", x"03", x"01", x"0a", x"fd", x"00",
    x"06", x"fc", x"08", x"05", x"23", x"3b", x"2c", x"e8",
    x"d0", x"dc", x"e4", x"e3", x"22", x"f4", x"df", x"ff",
    x"ea", x"cb", x"df", x"2e", x"f7", x"ec", x"05", x"cb",
    x"e2", x"05", x"1a", x"32", x"42", x"2c", x"2e", x"f9",
    x"0c", x"24", x"2a", x"0c", x"0b", x"bf", x"91", x"a3",
    x"0a", x"f5", x"05", x"2c", x"28", x"31", x"2f", x"f2",
    x"06", x"32", x"27", x"18", x"27", x"17", x"0b", x"15",
    x"12", x"24", x"fa", x"4b", x"38", x"25", x"24", x"2b",
    x"ab", x"e4", x"d5", x"f6", x"07", x"34", x"09", x"0d",
    x"d4", x"da", x"e5", x"0b", x"05", x"00", x"07", x"0e",
    x"fc", x"fe", x"06", x"02", x"fd", x"c8", x"db", x"c9",
    x"0e", x"08", x"ed", x"13", x"13", x"fd", x"13", x"bb",
    x"d9", x"2e", x"fa", x"d8", x"56", x"18", x"fb", x"2f",
    x"fa", x"13", x"0d", x"0e", x"13", x"19", x"10", x"2c",
    x"fc", x"ff", x"fc", x"ff", x"ff", x"fe", x"05", x"02",
    x"ff", x"08", x"ee", x"03", x"12", x"16", x"33", x"43",
    x"1a", x"37", x"d6", x"7d", x"ed", x"ef", x"a4", x"93",
    x"d1", x"e2", x"db", x"3a", x"bc", x"7f", x"5a", x"d7",
    x"ec", x"42", x"1b", x"3c", x"b3", x"c8", x"bc", x"24",
    x"0b", x"1b", x"fd", x"0e", x"19", x"aa", x"a4", x"a7",
    x"d7", x"bd", x"b2", x"e4", x"03", x"2d", x"bf", x"a2",
    x"0e", x"0d", x"00", x"2c", x"1f", x"10", x"d8", x"07",
    x"23", x"05", x"2e", x"2e", x"1b", x"31", x"31", x"11",
    x"f8", x"04", x"fe", x"04", x"06", x"00", x"fc", x"fe",
    x"04", x"fd", x"01", x"ff", x"fb", x"02", x"fe", x"01",
    x"fc", x"ff", x"44", x"3a", x"1a", x"f9", x"2b", x"2f",
    x"fc", x"f7", x"0c", x"ed", x"f8", x"db", x"03", x"25",
    x"28", x"f7", x"18", x"41", x"0b", x"03", x"17", x"11",
    x"15", x"3a", x"d6", x"0f", x"f5", x"11", x"20", x"01",
    x"f2", x"10", x"1c", x"63", x"81", x"d8", x"36", x"12",
    x"1c", x"22", x"2a", x"0c", x"f7", x"18", x"0a", x"c0",
    x"ad", x"fe", x"f3", x"f9", x"cf", x"2f", x"cf", x"fa",
    x"1b", x"d6", x"25", x"c6", x"bb", x"c2", x"63", x"ed",
    x"f2", x"15", x"16", x"19", x"f3", x"ef", x"e1", x"0a",
    x"e5", x"e0", x"f7", x"39", x"57", x"f1", x"31", x"4f",
    x"3f", x"ee", x"e2", x"3e", x"0a", x"00", x"39", x"1a",
    x"17", x"a1", x"d0", x"d9", x"19", x"09", x"e0", x"ca",
    x"a5", x"af", x"ef", x"ad", x"a8", x"dc", x"ed", x"16",
    x"d9", x"ee", x"11", x"cb", x"28", x"42", x"33", x"16",
    x"08", x"0a", x"18", x"2c", x"f3", x"fb", x"01", x"ef",
    x"3b", x"40", x"c4", x"10", x"2f", x"cd", x"9b", x"11",
    x"fb", x"fd", x"03", x"f7", x"fc", x"fd", x"f7", x"ff",
    x"fc", x"02", x"fa", x"fb", x"01", x"00", x"f9", x"fd",
    x"02", x"01", x"05", x"fe", x"fd", x"f8", x"01", x"fd",
    x"f7", x"fd", x"fb", x"fd", x"f6", x"fc", x"ff", x"fd",
    x"fd", x"f5", x"fa", x"fc", x"ff", x"00", x"fe", x"02",
    x"ff", x"fb", x"01", x"f8", x"fb", x"00", x"01", x"ff",
    x"03", x"00", x"08", x"04", x"fb", x"fb", x"fc", x"fc",
    x"fd", x"02", x"fb", x"fc", x"fe", x"fd", x"f7", x"ff",
    x"04", x"00", x"00", x"05", x"03", x"f8", x"fa", x"fb",
    x"fc", x"fe", x"fd", x"fc", x"ff", x"03", x"00", x"f9",
    x"02", x"f8", x"f5", x"f9", x"fc", x"00", x"03", x"01",
    x"fd", x"fe", x"05", x"fc", x"01", x"fd", x"04", x"fa",
    x"02", x"00", x"00", x"fc", x"01", x"fd", x"fd", x"01",
    x"f7", x"00", x"01", x"fd", x"00", x"fe", x"fc", x"fd",
    x"01", x"fa", x"fd", x"f9", x"f8", x"fe", x"fd", x"01",
    x"fe", x"00", x"01", x"fb", x"ff", x"00", x"fe", x"03",
    x"01", x"fb", x"02", x"fc", x"00", x"fa", x"00", x"ff",
    x"00", x"fa", x"fa", x"fe", x"fe", x"00", x"fc", x"ff",
    x"fc", x"fe", x"fc", x"fc", x"fc", x"01", x"fe", x"01",
    x"fb", x"00", x"04", x"fc", x"01", x"ff", x"ff", x"fb",
    x"fc", x"fb", x"02", x"03", x"ff", x"fe", x"03", x"01",
    x"fb", x"fb", x"ff", x"fc", x"fc", x"fe", x"fd", x"f9",
    x"01", x"0a", x"08", x"fe", x"fc", x"f6", x"fd", x"fe",
    x"fc", x"fc", x"fa", x"00", x"f8", x"fb", x"01", x"fc",
    x"fb", x"f7", x"00", x"02", x"02", x"fd", x"fd", x"ff",
    x"fe", x"f9", x"ff", x"fe", x"fe", x"01", x"03", x"00",
    x"ff", x"f9", x"fc", x"01", x"f7", x"fb", x"00", x"fe",
    x"05", x"03", x"f9", x"00", x"03", x"f7", x"02", x"01",
    x"fc", x"ff", x"00", x"f7", x"ff", x"02", x"ff", x"05",
    x"ff", x"f8", x"fb", x"fa", x"fd", x"00", x"fa", x"02",
    x"02", x"ff", x"fb", x"02", x"04", x"03", x"03", x"fe",
    x"02", x"fd", x"fc", x"02", x"01", x"fb", x"00", x"fd",
    x"01", x"fe", x"fd", x"f8", x"f9", x"fc", x"fb", x"f9",
    x"fe", x"fe", x"fc", x"01", x"fc", x"fe", x"00", x"fc",
    x"fa", x"fa", x"00", x"fd", x"00", x"ff", x"01", x"fc",
    x"fd", x"fb", x"fa", x"01", x"f9", x"f8", x"fc", x"00",
    x"00", x"f9", x"01", x"fa", x"f9", x"ff", x"fd", x"fd",
    x"fe", x"f8", x"f9", x"ff", x"fc", x"0b", x"fa", x"01",
    x"00", x"05", x"fd", x"03", x"01", x"fb", x"ff", x"00",
    x"fb", x"f8", x"02", x"f9", x"fd", x"fa", x"00", x"fa",
    x"ff", x"ff", x"02", x"fd", x"01", x"01", x"fe", x"00",
    x"ff", x"fb", x"03", x"fe", x"00", x"ff", x"fa", x"02",
    x"fe", x"f8", x"f7", x"fc", x"fc", x"ff", x"fd", x"00",
    x"00", x"ff", x"fa", x"fb", x"ff", x"00", x"fc", x"f5",
    x"01", x"f7", x"ff", x"fe", x"01", x"fa", x"fa", x"fd",
    x"fd", x"fb", x"01", x"01", x"fb", x"00", x"fd", x"01",
    x"00", x"03", x"fd", x"fe", x"fe", x"00", x"00", x"fe",
    x"fe", x"fb", x"03", x"fc", x"fc", x"fd", x"ff", x"fb",
    x"01", x"ff", x"f7", x"02", x"fd", x"fd", x"fb", x"02",
    x"f9", x"fc", x"fc", x"ff", x"ff", x"fe", x"01", x"fb",
    x"01", x"fa", x"fd", x"fc", x"02", x"01", x"fb", x"fd",
    x"03", x"fb", x"04", x"f7", x"f7", x"fe", x"01", x"fe",
    x"02", x"00", x"05", x"fb", x"03", x"fe", x"fd", x"03",
    x"01", x"ff", x"03", x"ff", x"01", x"fb", x"f9", x"00",
    x"fd", x"01", x"ff", x"03", x"00", x"03", x"03", x"fd",
    x"fd", x"05", x"fd", x"fb", x"fe", x"03", x"04", x"fe",
    x"02", x"04", x"01", x"00", x"03", x"00", x"ff", x"00",
    x"fd", x"ff", x"fd", x"00", x"f8", x"03", x"f9", x"01",
    x"fe", x"f7", x"f9", x"06", x"fd", x"fc", x"fc", x"f6",
    x"01", x"06", x"fd", x"ff", x"02", x"01", x"f6", x"fa",
    x"fd", x"f9", x"fc", x"01", x"fc", x"fd", x"00", x"fc",
    x"00", x"04", x"fa", x"04", x"fb", x"00", x"fd", x"ff",
    x"02", x"f9", x"fe", x"fe", x"f9", x"04", x"04", x"f9",
    x"00", x"fe", x"fc", x"f9", x"05", x"f9", x"01", x"fd",
    x"02", x"02", x"fd", x"fe", x"f7", x"fd", x"fc", x"00",
    x"f8", x"fe", x"03", x"01", x"f7", x"fd", x"fd", x"09",
    x"f9", x"fc", x"ff", x"fe", x"f7", x"fc", x"f8", x"ff",
    x"fb", x"fa", x"fd", x"f8", x"01", x"fb", x"f9", x"05",
    x"04", x"f8", x"fb", x"02", x"ff", x"05", x"fe", x"f8",
    x"01", x"fe", x"fc", x"ff", x"fa", x"fe", x"fd", x"04",
    x"fe", x"03", x"fe", x"f6", x"00", x"f8", x"fa", x"03",
    x"02", x"fd", x"01", x"f9", x"fa", x"ff", x"fe", x"06",
    x"04", x"fc", x"02", x"fb", x"fe", x"fb", x"04", x"00",
    x"03", x"04", x"ff", x"02", x"07", x"fa", x"fb", x"fe",
    x"04", x"fb", x"02", x"00", x"04", x"ff", x"01", x"fc",
    x"fe", x"03", x"fa", x"f6", x"fd", x"ff", x"fd", x"01",
    x"f8", x"fa", x"fc", x"fe", x"03", x"00", x"03", x"02",
    x"fb", x"fb", x"ff", x"03", x"fe", x"02", x"fb", x"fd",
    x"00", x"fb", x"ff", x"05", x"ff", x"02", x"fb", x"fa",
    x"fc", x"fc", x"fe", x"04", x"fc", x"ff", x"ff", x"fa",
    x"fe", x"fa", x"fa", x"03", x"fa", x"fc", x"fa", x"fb",
    x"02", x"03", x"02", x"01", x"fd", x"fe", x"fc", x"fc",
    x"00", x"ff", x"00", x"ff", x"fa", x"fa", x"01", x"03",
    x"ff", x"fe", x"fb", x"01", x"f9", x"fe", x"07", x"fa",
    x"02", x"fb", x"fc", x"fc", x"ff", x"00", x"01", x"03",
    x"04", x"ff", x"fd", x"02", x"04", x"fc", x"04", x"fa",
    x"fa", x"ff", x"fe", x"fe", x"03", x"ff", x"02", x"03",
    x"04", x"03", x"01", x"03", x"fe", x"fb", x"fd", x"01",
    x"fd", x"fd", x"fd", x"04", x"fb", x"fb", x"fd", x"fd",
    x"01", x"01", x"04", x"02", x"03", x"04", x"01", x"02",
    x"00", x"fe", x"fd", x"ff", x"fe", x"fd", x"fc", x"01",
    x"fd", x"fc", x"03", x"fe", x"fd", x"ff", x"02", x"01",
    x"fe", x"03", x"fe", x"fc", x"fd", x"02", x"02", x"fb",
    x"fe", x"fc", x"fa", x"ff", x"fa", x"fd", x"04", x"fe",
    x"03", x"fb", x"fc", x"00", x"fc", x"fa", x"fe", x"fc",
    x"ff", x"fb", x"fd", x"04", x"fa", x"00", x"fe", x"fc",
    x"04", x"01", x"fa", x"ff", x"fa", x"f8", x"fd", x"fc",
    x"03", x"fe", x"01", x"fe", x"00", x"ff", x"fe", x"fa",
    x"fe", x"fc", x"fa", x"fa", x"fc", x"06", x"03", x"f8",
    x"00", x"ff", x"02", x"fe", x"fe", x"00", x"01", x"fe",
    x"fd", x"00", x"02", x"fc", x"00", x"03", x"00", x"01",
    x"fc", x"fe", x"fb", x"fb", x"01", x"fe", x"fe", x"fc",
    x"04", x"fa", x"fa", x"fc", x"fb", x"fe", x"fd", x"fd",
    x"00", x"04", x"04", x"03", x"00", x"03", x"fd", x"02",
    x"ff", x"fb", x"ff", x"fb", x"fa", x"fb", x"04", x"fa",
    x"02", x"fc", x"ff", x"fe", x"01", x"ff", x"fa", x"03",
    x"00", x"01", x"00", x"04", x"ff", x"ff", x"01", x"fc",
    x"01", x"fe", x"03", x"fe", x"fc", x"ff", x"fd", x"fe",
    x"fb", x"fd", x"fe", x"fa", x"fe", x"00", x"01", x"00",
    x"f6", x"fa", x"fb", x"ff", x"fd", x"fd", x"fe", x"01",
    x"fd", x"ff", x"fa", x"ff", x"fb", x"01", x"04", x"fb",
    x"01", x"fe", x"fb", x"fb", x"ff", x"fd", x"01", x"fe",
    x"fc", x"fa", x"01", x"fd", x"03", x"fe", x"fb", x"fb",
    x"fe", x"01", x"01", x"05", x"03", x"01", x"fe", x"01",
    x"02", x"02", x"02", x"fc", x"01", x"fd", x"03", x"ff",
    x"03", x"fb", x"02", x"fa", x"fe", x"fd", x"fc", x"00",
    x"03", x"00", x"fc", x"fa", x"fd", x"fc", x"fc", x"fd",
    x"fd", x"00", x"fd", x"fc", x"04", x"fe", x"fb", x"04",
    x"04", x"ff", x"00", x"04", x"03", x"fb", x"fa", x"00",
    x"fa", x"00", x"fb", x"01", x"01", x"fb", x"02", x"00",
    x"fd", x"fb", x"00", x"fe", x"fc", x"fb", x"fe", x"fb",
    x"04", x"fd", x"fa", x"ff", x"01", x"fc", x"ff", x"00",
    x"fa", x"fe", x"fb", x"04", x"00", x"05", x"fa", x"ff",
    x"00", x"fe", x"01", x"fa", x"fa", x"02", x"fb", x"ff",
    x"01", x"02", x"01", x"ff", x"fc", x"04", x"01", x"fa",
    x"03", x"04", x"00", x"fb", x"fd", x"06", x"ff", x"02",
    x"00", x"fb", x"00", x"03", x"01", x"fc", x"04", x"01",
    x"ff", x"fe", x"01", x"fc", x"02", x"02", x"ff", x"00",
    x"03", x"fc", x"03", x"02", x"fd", x"04", x"02", x"03",
    x"ff", x"fc", x"ff", x"fb", x"fc", x"00", x"fb", x"03",
    x"01", x"fd", x"02", x"f9", x"01", x"fd", x"02", x"00",
    x"ff", x"fa", x"fd", x"ff", x"fe", x"fc", x"fd", x"01",
    x"01", x"fd", x"fe", x"03", x"fb", x"00", x"fe", x"fe",
    x"03", x"fc", x"fa", x"fb", x"02", x"03", x"01", x"01",
    x"fd", x"02", x"fd", x"01", x"01", x"01", x"fc", x"fe",
    x"00", x"04", x"ff", x"fb", x"04", x"ff", x"ff", x"fb",
    x"fb", x"fb", x"fb", x"ff", x"fe", x"ff", x"ff", x"02",
    x"ff", x"00", x"fe", x"fd", x"02", x"fa", x"02", x"fd",
    x"fe", x"00", x"fa", x"fc", x"fa", x"01", x"fb", x"fc",
    x"f9", x"05", x"ff", x"fe", x"fb", x"fd", x"fb", x"00",
    x"03", x"fb", x"fd", x"fe", x"04", x"fd", x"fd", x"fa",
    x"ff", x"fd", x"fb", x"fa", x"03", x"f9", x"fe", x"fd",
    x"fa", x"04", x"fe", x"00", x"fb", x"ff", x"fc", x"fe",
    x"fb", x"ff", x"ff", x"04", x"01", x"01", x"ff", x"fe",
    x"1f", x"fb", x"f8", x"0d", x"00", x"1f", x"c5", x"ce",
    x"23", x"f7", x"18", x"11", x"0d", x"ec", x"f8", x"f8",
    x"cb", x"bf", x"db", x"e3", x"ef", x"e3", x"e5", x"ff",
    x"ce", x"db", x"1a", x"d6", x"e9", x"d8", x"aa", x"ea",
    x"fd", x"3b", x"18", x"0e", x"21", x"2e", x"1f", x"09",
    x"0d", x"21", x"d4", x"cc", x"ae", x"f8", x"0d", x"e2",
    x"19", x"e2", x"e1", x"1d", x"f5", x"e9", x"d4", x"0a",
    x"19", x"08", x"01", x"d0", x"f5", x"f9", x"24", x"a8",
    x"ac", x"1c", x"04", x"01", x"3c", x"24", x"1b", x"f3",
    x"c1", x"bf", x"b9", x"f0", x"02", x"3b", x"ea", x"1f",
    x"0a", x"18", x"07", x"cd", x"d7", x"c5", x"ed", x"14",
    x"ee", x"cf", x"fa", x"f3", x"ce", x"83", x"2d", x"11",
    x"24", x"16", x"3e", x"4c", x"38", x"db", x"18", x"39",
    x"fc", x"3e", x"63", x"16", x"f9", x"f8", x"24", x"02",
    x"e0", x"e1", x"dd", x"d9", x"f2", x"c0", x"5f", x"19",
    x"f9", x"f7", x"d6", x"13", x"36", x"1f", x"df", x"d2",
    x"bf", x"b9", x"e8", x"f2", x"ea", x"1d", x"26", x"ed",
    x"1f", x"e9", x"e6", x"da", x"f0", x"a3", x"a8", x"b7",
    x"f2", x"01", x"01", x"fc", x"f3", x"d5", x"03", x"24",
    x"4e", x"fb", x"ff", x"04", x"04", x"fc", x"03", x"03",
    x"01", x"03", x"0c", x"31", x"db", x"08", x"2b", x"c0",
    x"21", x"3d", x"16", x"03", x"10", x"1c", x"06", x"ff",
    x"1a", x"20", x"f4", x"d9", x"db", x"f1", x"91", x"15",
    x"e2", x"be", x"26", x"f6", x"d1", x"f6", x"03", x"08",
    x"ee", x"1a", x"25", x"b1", x"e3", x"2d", x"f6", x"03",
    x"01", x"e9", x"f1", x"23", x"ac", x"a7", x"16", x"2e",
    x"18", x"d9", x"20", x"32", x"2c", x"fc", x"e1", x"ed",
    x"5e", x"0e", x"fa", x"23", x"d6", x"17", x"18", x"17",
    x"35", x"d2", x"e2", x"af", x"fb", x"ea", x"0d", x"22",
    x"01", x"27", x"e0", x"f3", x"ee", x"18", x"31", x"1b",
    x"b9", x"c8", x"e8", x"f9", x"fd", x"fd", x"fe", x"00",
    x"00", x"ff", x"00", x"02", x"f0", x"97", x"ce", x"0f",
    x"f8", x"fe", x"06", x"ff", x"19", x"36", x"1d", x"0e",
    x"15", x"21", x"0a", x"1d", x"ee", x"d4", x"14", x"0b",
    x"c6", x"ee", x"d6", x"e1", x"38", x"13", x"f5", x"fe",
    x"03", x"15", x"eb", x"ec", x"df", x"10", x"25", x"f9",
    x"ed", x"2d", x"de", x"28", x"1e", x"5c", x"fa", x"39",
    x"7a", x"10", x"ef", x"14", x"0d", x"d3", x"db", x"0d",
    x"0c", x"e2", x"22", x"e6", x"08", x"38", x"04", x"26",
    x"35", x"49", x"4c", x"0a", x"b0", x"ee", x"04", x"d6",
    x"f9", x"f9", x"b2", x"c8", x"02", x"ff", x"fd", x"08",
    x"14", x"f8", x"03", x"0e", x"fc", x"ff", x"e8", x"dd",
    x"0b", x"f6", x"f4", x"14", x"ea", x"eb", x"d4", x"e5",
    x"c5", x"d8", x"17", x"f3", x"65", x"41", x"5c", x"a9",
    x"ee", x"08", x"f6", x"e4", x"bf", x"6d", x"47", x"48",
    x"fb", x"05", x"ff", x"fc", x"00", x"ff", x"02", x"fb",
    x"04", x"22", x"ca", x"da", x"12", x"0f", x"01", x"15",
    x"e6", x"f8", x"e7", x"b7", x"9f", x"ea", x"ff", x"05",
    x"1e", x"32", x"41", x"0e", x"f2", x"03", x"33", x"20",
    x"15", x"dd", x"f2", x"fd", x"a9", x"b2", x"e0", x"f7",
    x"e7", x"e1", x"1d", x"ee", x"fa", x"ee", x"e8", x"1a",
    x"2d", x"0d", x"0c", x"1b", x"01", x"21", x"f3", x"ba",
    x"f4", x"d8", x"f7", x"ba", x"ee", x"dc", x"d9", x"1e",
    x"14", x"27", x"21", x"01", x"13", x"20", x"f5", x"19",
    x"fb", x"01", x"07", x"01", x"fe", x"04", x"f9", x"0a",
    x"04", x"fc", x"02", x"fe", x"fb", x"00", x"04", x"ff",
    x"07", x"fd", x"e5", x"b2", x"b4", x"1c", x"fa", x"f7",
    x"bd", x"ba", x"bb", x"d2", x"47", x"d1", x"1f", x"1a",
    x"20", x"24", x"59", x"69", x"39", x"04", x"d3", x"14",
    x"01", x"0b", x"fd", x"2c", x"e2", x"0d", x"06", x"0b",
    x"10", x"22", x"2f", x"f0", x"0f", x"e4", x"d9", x"bd",
    x"f9", x"e4", x"36", x"3d", x"20", x"3d", x"0b", x"48",
    x"2d", x"27", x"1c", x"09", x"ef", x"e8", x"f3", x"f4",
    x"31", x"1a", x"12", x"27", x"06", x"04", x"f6", x"25",
    x"1c", x"0d", x"df", x"fa", x"1f", x"fd", x"f3", x"1e",
    x"0a", x"c4", x"ce", x"db", x"f2", x"d9", x"be", x"eb",
    x"f1", x"a7", x"ea", x"0e", x"14", x"11", x"bd", x"ed",
    x"e4", x"3d", x"19", x"ec", x"3b", x"e3", x"df", x"39",
    x"1c", x"18", x"f3", x"c7", x"c1", x"04", x"0e", x"c2",
    x"dd", x"ff", x"e2", x"dc", x"ce", x"ec", x"c4", x"eb",
    x"11", x"00", x"e3", x"f1", x"0f", x"ed", x"d4", x"44",
    x"3d", x"52", x"11", x"e3", x"0f", x"34", x"0d", x"25",
    x"ec", x"f4", x"ca", x"23", x"06", x"03", x"f7", x"b5",
    x"04", x"02", x"dd", x"c2", x"f3", x"11", x"28", x"cb",
    x"f1", x"ec", x"f3", x"eb", x"a5", x"d2", x"c4", x"e9",
    x"dc", x"e0", x"ec", x"0a", x"02", x"05", x"da", x"c4",
    x"eb", x"ce", x"d6", x"ef", x"aa", x"cd", x"00", x"04",
    x"2f", x"26", x"8c", x"a1", x"bc", x"b5", x"15", x"10",
    x"d8", x"fa", x"11", x"d1", x"06", x"1d", x"e8", x"03",
    x"11", x"09", x"04", x"f5", x"c5", x"f1", x"19", x"c5",
    x"f7", x"dc", x"41", x"4c", x"58", x"3e", x"4b", x"0f",
    x"b5", x"fc", x"0d", x"f8", x"fc", x"10", x"fd", x"00",
    x"ef", x"06", x"24", x"3e", x"08", x"06", x"f5", x"22",
    x"1f", x"d7", x"f9", x"f1", x"f7", x"36", x"e7", x"c6",
    x"37", x"f2", x"e5", x"1f", x"da", x"da", x"42", x"fb",
    x"f9", x"2d", x"d8", x"f6", x"1a", x"f6", x"26", x"1b",
    x"e9", x"ec", x"e4", x"bc", x"d2", x"ad", x"44", x"6a",
    x"d8", x"c6", x"9d", x"2b", x"0a", x"d8", x"a6", x"8b",
    x"89", x"9f", x"99", x"ba", x"4a", x"42", x"0a", x"c2",
    x"45", x"27", x"00", x"21", x"11", x"d3", x"cf", x"e3",
    x"2a", x"20", x"f7", x"f9", x"1b", x"18", x"ee", x"03",
    x"ff", x"05", x"fe", x"fe", x"05", x"05", x"ff", x"05",
    x"01", x"01", x"92", x"9d", x"22", x"e4", x"ec", x"c9",
    x"47", x"41", x"2a", x"06", x"e0", x"fd", x"00", x"fd",
    x"12", x"54", x"16", x"33", x"ed", x"ea", x"c9", x"de",
    x"c8", x"a2", x"24", x"ec", x"0e", x"e5", x"dd", x"e8",
    x"f1", x"f9", x"ef", x"10", x"1c", x"24", x"d7", x"fc",
    x"dc", x"00", x"ea", x"e8", x"e1", x"fb", x"14", x"ee",
    x"f0", x"b9", x"f3", x"2f", x"df", x"20", x"18", x"e3",
    x"d8", x"d4", x"c9", x"4d", x"0f", x"12", x"2d", x"29",
    x"2a", x"0f", x"e9", x"cb", x"f4", x"11", x"f6", x"10",
    x"ee", x"2c", x"d2", x"e9", x"05", x"01", x"0a", x"06",
    x"10", x"4f", x"21", x"00", x"02", x"ff", x"f8", x"fa",
    x"fd", x"ff", x"ff", x"f7", x"ed", x"1a", x"cc", x"03",
    x"0b", x"e6", x"1e", x"3a", x"13", x"f6", x"d5", x"e1",
    x"11", x"12", x"d5", x"00", x"e7", x"a9", x"fb", x"b6",
    x"91", x"de", x"e4", x"b5", x"1c", x"17", x"1b", x"ca",
    x"d5", x"f6", x"f8", x"f6", x"14", x"fc", x"07", x"18",
    x"bc", x"95", x"e6", x"2c", x"28", x"f5", x"0f", x"2c",
    x"58", x"17", x"05", x"f9", x"1d", x"0d", x"32", x"0f",
    x"22", x"98", x"b5", x"da", x"ec", x"2d", x"1a", x"10",
    x"2e", x"03", x"fe", x"b8", x"02", x"0f", x"32", x"2e",
    x"e3", x"1e", x"13", x"e7", x"f9", x"01", x"ff", x"fa",
    x"ff", x"01", x"02", x"03", x"08", x"c4", x"a1", x"a3",
    x"0a", x"ec", x"00", x"e1", x"f4", x"18", x"22", x"0f",
    x"f4", x"1f", x"d5", x"d6", x"aa", x"1e", x"42", x"e0",
    x"13", x"34", x"12", x"bf", x"d9", x"bf", x"01", x"20",
    x"fd", x"01", x"02", x"03", x"00", x"fc", x"02", x"ff",
    x"fb", x"45", x"d6", x"95", x"a4", x"aa", x"c5", x"fa",
    x"ff", x"05", x"a5", x"89", x"cf", x"05", x"df", x"e9",
    x"2c", x"24", x"11", x"02", x"d9", x"d7", x"2d", x"07",
    x"07", x"46", x"1d", x"e9", x"ed", x"d2", x"c8", x"e3",
    x"dc", x"ec", x"20", x"03", x"08", x"c0", x"b9", x"b6",
    x"f9", x"f9", x"f6", x"27", x"0c", x"0f", x"d3", x"03",
    x"1c", x"00", x"e9", x"11", x"02", x"da", x"af", x"db",
    x"12", x"1f", x"f0", x"13", x"f8", x"3d", x"22", x"26",
    x"fd", x"00", x"05", x"02", x"06", x"03", x"03", x"02",
    x"01", x"fe", x"09", x"05", x"03", x"04", x"07", x"03",
    x"f8", x"03", x"f6", x"2d", x"27", x"ee", x"26", x"26",
    x"ca", x"c9", x"cd", x"ad", x"c8", x"c0", x"db", x"18",
    x"ce", x"1e", x"58", x"9a", x"c8", x"fe", x"09", x"fc",
    x"1a", x"07", x"f8", x"14", x"e9", x"e6", x"12", x"ec",
    x"27", x"02", x"19", x"08", x"1b", x"07", x"80", x"e2",
    x"ed", x"29", x"e8", x"e1", x"40", x"14", x"cf", x"f6",
    x"ea", x"de", x"2f", x"1d", x"e1", x"df", x"f6", x"f4",
    x"e1", x"f8", x"cf", x"11", x"01", x"dc", x"02", x"d3",
    x"d8", x"65", x"f6", x"fe", x"29", x"29", x"24", x"cf",
    x"c1", x"c7", x"e0", x"25", x"ff", x"c6", x"ef", x"06",
    x"cd", x"c4", x"1e", x"ed", x"1b", x"23", x"e9", x"f0",
    x"ed", x"18", x"18", x"f5", x"da", x"3b", x"3c", x"07",
    x"53", x"40", x"13", x"ea", x"87", x"de", x"07", x"f1",
    x"27", x"17", x"03", x"07", x"e3", x"b4", x"e5", x"e8",
    x"b0", x"09", x"f8", x"08", x"fa", x"f2", x"f8", x"bf",
    x"dc", x"d1", x"1c", x"15", x"08", x"07", x"13", x"2c",
    x"ef", x"03", x"20", x"bf", x"d0", x"17", x"34", x"4b",
    x"5c", x"17", x"23", x"22", x"de", x"ef", x"fc", x"e4",
    x"27", x"28", x"23", x"f5", x"d3", x"c7", x"17", x"45",
    x"49", x"48", x"53", x"ee", x"d4", x"03", x"17", x"01",
    x"21", x"d7", x"c1", x"e7", x"eb", x"e7", x"f8", x"e6",
    x"f5", x"22", x"1e", x"3c", x"61", x"15", x"2d", x"0d",
    x"26", x"ee", x"b7", x"c6", x"fe", x"0b", x"2f", x"28",
    x"3b", x"ec", x"2c", x"23", x"f6", x"dd", x"d4", x"e1",
    x"f1", x"66", x"ca", x"d3", x"ac", x"98", x"b4", x"1a",
    x"e6", x"08", x"db", x"16", x"08", x"e9", x"ff", x"12",
    x"22", x"1c", x"02", x"1b", x"38", x"34", x"f6", x"d3",
    x"f8", x"e3", x"24", x"29", x"31", x"3b", x"33", x"10",
    x"4e", x"4d", x"4a", x"e9", x"fe", x"1f", x"f4", x"fd",
    x"2e", x"ea", x"f0", x"eb", x"e4", x"f7", x"f8", x"dd",
    x"15", x"21", x"ce", x"04", x"25", x"d5", x"e3", x"e1",
    x"1e", x"28", x"f0", x"15", x"1f", x"f3", x"21", x"f3",
    x"37", x"d7", x"b9", x"d1", x"dd", x"b8", x"d3", x"e3",
    x"de", x"f1", x"05", x"17", x"0c", x"2f", x"1a", x"ea",
    x"f5", x"16", x"d0", x"10", x"ed", x"ab", x"0b", x"d8",
    x"e2", x"00", x"01", x"fc", x"06", x"fc", x"05", x"03",
    x"05", x"fe", x"2d", x"62", x"1d", x"f2", x"08", x"ba",
    x"a6", x"64", x"bb", x"00", x"f4", x"15", x"17", x"23",
    x"16", x"01", x"0a", x"cf", x"06", x"07", x"2c", x"16",
    x"22", x"09", x"f4", x"f6", x"df", x"db", x"0d", x"1d",
    x"00", x"10", x"04", x"03", x"03", x"16", x"f0", x"0e",
    x"1d", x"13", x"ed", x"d4", x"1b", x"3d", x"44", x"fc",
    x"e1", x"f6", x"f7", x"ec", x"05", x"25", x"25", x"27",
    x"cf", x"9b", x"d8", x"ba", x"d0", x"f0", x"d7", x"73",
    x"38", x"f0", x"03", x"04", x"02", x"01", x"14", x"fe",
    x"fd", x"f4", x"0d", x"e9", x"00", x"0c", x"16", x"07",
    x"29", x"1b", x"1d", x"00", x"fd", x"02", x"03", x"00",
    x"ff", x"03", x"03", x"01", x"0d", x"15", x"03", x"f3",
    x"e7", x"d8", x"dc", x"f3", x"f0", x"07", x"18", x"33",
    x"1c", x"3b", x"ee", x"40", x"03", x"b0", x"f5", x"03",
    x"dd", x"0f", x"0f", x"19", x"e7", x"dd", x"f8", x"cf",
    x"b9", x"f3", x"18", x"06", x"02", x"d1", x"e7", x"dd",
    x"0e", x"5b", x"3a", x"0e", x"1c", x"2c", x"ce", x"dd",
    x"16", x"d6", x"00", x"ef", x"15", x"0d", x"ff", x"f1",
    x"de", x"f8", x"08", x"f9", x"45", x"ee", x"de", x"f9",
    x"c0", x"c1", x"08", x"0a", x"ef", x"e4", x"e1", x"02",
    x"f0", x"3f", x"ea", x"f5", x"f4", x"f7", x"fb", x"f9",
    x"ec", x"01", x"f1", x"f3", x"fe", x"e9", x"0f", x"47",
    x"1e", x"05", x"19", x"1e", x"eb", x"ae", x"3b", x"d4",
    x"bc", x"13", x"1d", x"14", x"1c", x"33", x"0e", x"21",
    x"56", x"56", x"be", x"f7", x"f8", x"18", x"fa", x"e4",
    x"fc", x"01", x"fc", x"ff", x"03", x"fe", x"fe", x"07",
    x"01", x"e4", x"f0", x"f8", x"d3", x"12", x"31", x"0b",
    x"df", x"dc", x"34", x"c0", x"a7", x"cd", x"e4", x"15",
    x"f2", x"11", x"0f", x"fe", x"21", x"0c", x"29", x"e9",
    x"df", x"34", x"f6", x"04", x"05", x"ff", x"62", x"28",
    x"45", x"60", x"16", x"1f", x"ee", x"b3", x"b3", x"ea",
    x"f7", x"29", x"57", x"0e", x"1e", x"55", x"3a", x"23",
    x"ed", x"e9", x"c2", x"ae", x"04", x"c7", x"de", x"28",
    x"52", x"39", x"0d", x"24", x"fb", x"f2", x"fa", x"30",
    x"01", x"fb", x"fe", x"01", x"00", x"00", x"fd", x"00",
    x"07", x"03", x"02", x"0b", x"05", x"fe", x"ff", x"02",
    x"02", x"fd", x"1c", x"19", x"28", x"e3", x"8c", x"b4",
    x"1a", x"41", x"1d", x"e9", x"4a", x"f5", x"01", x"fd",
    x"13", x"d4", x"03", x"c8", x"1e", x"2e", x"25", x"1b",
    x"36", x"15", x"d0", x"e6", x"c1", x"f0", x"eb", x"01",
    x"bc", x"f1", x"10", x"34", x"27", x"0e", x"01", x"54",
    x"3e", x"f6", x"24", x"2b", x"eb", x"04", x"eb", x"c6",
    x"ab", x"c6", x"14", x"2d", x"1f", x"13", x"da", x"e7",
    x"0f", x"00", x"2e", x"cc", x"e8", x"ff", x"fc", x"29",
    x"15", x"fb", x"f9", x"26", x"cc", x"c4", x"ea", x"f7",
    x"19", x"2d", x"dc", x"ef", x"3c", x"f9", x"ef", x"2a",
    x"1a", x"fc", x"fc", x"07", x"e0", x"1a", x"16", x"0e",
    x"dd", x"19", x"05", x"01", x"03", x"2e", x"d4", x"1c",
    x"6f", x"bc", x"0e", x"09", x"0b", x"2e", x"18", x"fb",
    x"dd", x"e5", x"c3", x"f2", x"e2", x"ff", x"e6", x"dc",
    x"ce", x"c2", x"b0", x"e1", x"ae", x"48", x"54", x"da",
    x"d8", x"c6", x"09", x"ea", x"e8", x"09", x"13", x"04",
    x"f8", x"c2", x"99", x"e4", x"bc", x"d9", x"f5", x"12",
    x"5b", x"07", x"0a", x"ef", x"a2", x"d3", x"f2", x"28",
    x"f5", x"e0", x"19", x"1d", x"0a", x"34", x"28", x"2c",
    x"0a", x"fe", x"2c", x"c5", x"ea", x"f1", x"f4", x"11",
    x"02", x"dd", x"f6", x"c6", x"15", x"03", x"03", x"01",
    x"09", x"ed", x"16", x"ec", x"07", x"31", x"d6", x"5b",
    x"2b", x"f7", x"de", x"9e", x"25", x"06", x"fe", x"f2",
    x"10", x"fa", x"ea", x"fa", x"28", x"24", x"1e", x"e6",
    x"1a", x"07", x"ab", x"be", x"0e", x"d2", x"fa", x"ec",
    x"da", x"f8", x"dc", x"f1", x"03", x"e2", x"17", x"2c",
    x"32", x"26", x"1a", x"02", x"c2", x"e8", x"06", x"fb",
    x"fe", x"0b", x"12", x"16", x"0a", x"6b", x"2b", x"24",
    x"29", x"04", x"09", x"cf", x"13", x"db", x"d3", x"03",
    x"08", x"08", x"07", x"ee", x"f8", x"13", x"e9", x"e2",
    x"b0", x"e8", x"14", x"e1", x"ec", x"15", x"ef", x"c1",
    x"2c", x"25", x"2d", x"20", x"30", x"48", x"44", x"29",
    x"2f", x"f9", x"f1", x"0c", x"04", x"17", x"08", x"1b",
    x"dc", x"e8", x"26", x"0b", x"e6", x"0f", x"08", x"f7",
    x"df", x"a5", x"b3", x"ca", x"dd", x"e1", x"f6", x"fb",
    x"f1", x"fc", x"03", x"03", x"fe", x"04", x"04", x"00",
    x"fd", x"00", x"25", x"0c", x"fd", x"22", x"00", x"f3",
    x"00", x"ef", x"06", x"10", x"0c", x"0a", x"0e", x"f0",
    x"ed", x"02", x"0a", x"0c", x"50", x"20", x"fe", x"1a",
    x"39", x"29", x"cb", x"2d", x"03", x"29", x"27", x"f2",
    x"1e", x"16", x"06", x"19", x"10", x"3c", x"f6", x"d3",
    x"df", x"27", x"ea", x"fc", x"e0", x"e8", x"f7", x"12",
    x"17", x"d2", x"22", x"f4", x"ea", x"dc", x"e5", x"f2",
    x"ce", x"b6", x"e6", x"d6", x"e6", x"0b", x"db", x"e7",
    x"1c", x"0b", x"10", x"29", x"07", x"03", x"00", x"32",
    x"2a", x"09", x"12", x"23", x"fd", x"15", x"14", x"16",
    x"f7", x"f9", x"24", x"fe", x"fe", x"fd", x"02", x"04",
    x"04", x"fb", x"00", x"fd", x"df", x"b4", x"e2", x"ff",
    x"bc", x"d4", x"cf", x"9f", x"c8", x"13", x"e1", x"b8",
    x"30", x"1e", x"ef", x"0a", x"06", x"05", x"3f", x"2e",
    x"0b", x"2b", x"16", x"3c", x"19", x"19", x"0a", x"a0",
    x"b7", x"b3", x"a4", x"7c", x"94", x"04", x"ca", x"e5",
    x"e6", x"18", x"f1", x"e2", x"ee", x"2e", x"e7", x"12",
    x"11", x"14", x"ec", x"fc", x"f8", x"05", x"bc", x"ef",
    x"f0", x"f8", x"e3", x"f3", x"0d", x"e0", x"13", x"18",
    x"2d", x"ea", x"fe", x"c1", x"b5", x"fa", x"b7", x"c8",
    x"f3", x"2f", x"47", x"26", x"08", x"07", x"0e", x"0a",
    x"07", x"10", x"03", x"03", x"02", x"48", x"38", x"19",
    x"40", x"fd", x"e4", x"0c", x"eb", x"e9", x"00", x"e6",
    x"c9", x"29", x"f7", x"cf", x"df", x"26", x"22", x"e6",
    x"dc", x"b2", x"02", x"f6", x"24", x"14", x"f8", x"1c",
    x"04", x"05", x"02", x"fe", x"fb", x"fd", x"05", x"04",
    x"03", x"14", x"02", x"23", x"33", x"23", x"1b", x"0b",
    x"2b", x"2a", x"bd", x"8f", x"a2", x"9c", x"8c", x"b3",
    x"c9", x"eb", x"05", x"71", x"15", x"1f", x"47", x"1d",
    x"1a", x"15", x"1b", x"2f", x"10", x"10", x"12", x"3e",
    x"16", x"0b", x"0c", x"0a", x"25", x"c5", x"c0", x"c1",
    x"a0", x"c9", x"f3", x"d6", x"02", x"3a", x"27", x"b5",
    x"bc", x"21", x"fb", x"ed", x"08", x"fd", x"dd", x"44",
    x"40", x"fb", x"2c", x"28", x"06", x"1d", x"31", x"4a",
    x"fc", x"fc", x"00", x"fe", x"03", x"04", x"04", x"fd",
    x"00", x"fc", x"02", x"fd", x"03", x"02", x"00", x"00",
    x"fd", x"fc", x"26", x"e9", x"d4", x"03", x"cb", x"be",
    x"fa", x"ce", x"f4", x"e6", x"ca", x"ca", x"0f", x"eb",
    x"04", x"25", x"26", x"0f", x"4a", x"56", x"30", x"30",
    x"25", x"24", x"dd", x"c8", x"e9", x"d7", x"ff", x"fd",
    x"11", x"05", x"04", x"f1", x"e8", x"00", x"1d", x"28",
    x"14", x"2b", x"04", x"e1", x"fa", x"03", x"fd", x"e2",
    x"a7", x"d7", x"66", x"fa", x"08", x"1e", x"0e", x"05",
    x"3a", x"dd", x"0c", x"00", x"f6", x"0c", x"f1", x"dd",
    x"e2", x"c5", x"1c", x"48", x"30", x"13", x"0d", x"3c",
    x"0a", x"e6", x"e5", x"f5", x"0f", x"2b", x"29", x"12",
    x"11", x"31", x"11", x"35", x"32", x"21", x"23", x"21",
    x"0a", x"c6", x"eb", x"eb", x"12", x"03", x"ff", x"f7",
    x"c5", x"cd", x"b6", x"ed", x"05", x"27", x"fb", x"d6",
    x"0b", x"1e", x"ea", x"d6", x"01", x"e2", x"d7", x"e5",
    x"13", x"8e", x"fa", x"18", x"db", x"01", x"2b", x"ae",
    x"ec", x"16", x"ef", x"be", x"be", x"03", x"d6", x"c0",
    x"09", x"2e", x"47", x"2c", x"22", x"06", x"da", x"ee",
    x"a5", x"e2", x"0b", x"19", x"44", x"0b", x"fc", x"3d",
    x"1a", x"ff", x"ff", x"30", x"25", x"05", x"2a", x"25",
    x"97", x"c4", x"e3", x"15", x"eb", x"de", x"dc", x"e2",
    x"d6", x"f0", x"da", x"03", x"f9", x"2c", x"3e", x"31",
    x"43", x"57", x"bf", x"c5", x"ba", x"fc", x"07", x"ed",
    x"ab", x"d1", x"c3", x"e5", x"fd", x"d0", x"e2", x"24",
    x"11", x"c5", x"c0", x"eb", x"f3", x"0e", x"0d", x"87",
    x"80", x"05", x"d9", x"b3", x"be", x"28", x"1f", x"00",
    x"25", x"03", x"11", x"d0", x"d6", x"01", x"f5", x"f0",
    x"f2", x"bb", x"d1", x"fa", x"02", x"e6", x"e5", x"d9",
    x"04", x"f6", x"22", x"f2", x"22", x"25", x"2e", x"f8",
    x"12", x"e4", x"d6", x"06", x"ee", x"06", x"ab", x"03",
    x"f7", x"b5", x"26", x"1a", x"36", x"2d", x"18", x"5b",
    x"2e", x"1a", x"c1", x"cd", x"e1", x"35", x"23", x"4e",
    x"f9", x"d7", x"e1", x"eb", x"0e", x"e1", x"15", x"d4",
    x"ca", x"db", x"bb", x"ce", x"cf", x"f3", x"e1", x"38",
    x"2e", x"37", x"26", x"2d", x"04", x"f8", x"19", x"0f",
    x"f3", x"de", x"d8", x"f6", x"e2", x"e8", x"46", x"3f",
    x"32", x"04", x"06", x"fd", x"04", x"00", x"ff", x"03",
    x"01", x"fd", x"c9", x"78", x"94", x"3d", x"14", x"8e",
    x"27", x"26", x"12", x"e1", x"ff", x"15", x"d7", x"e5",
    x"db", x"d5", x"be", x"df", x"14", x"0c", x"15", x"29",
    x"2d", x"fd", x"0d", x"0f", x"f5", x"df", x"09", x"16",
    x"bd", x"bb", x"93", x"02", x"d7", x"c1", x"8c", x"be",
    x"cc", x"20", x"0e", x"fb", x"66", x"43", x"20", x"3e",
    x"35", x"31", x"21", x"23", x"30", x"4e", x"2c", x"0f",
    x"af", x"06", x"ee", x"f7", x"40", x"13", x"0d", x"27",
    x"07", x"eb", x"ed", x"d2", x"fb", x"ec", x"09", x"b0",
    x"0e", x"28", x"cc", x"e4", x"ee", x"c3", x"93", x"80",
    x"05", x"cc", x"d6", x"00", x"01", x"01", x"00", x"05",
    x"04", x"ff", x"fc", x"03", x"42", x"f4", x"0e", x"d6",
    x"12", x"13", x"18", x"ff", x"f5", x"c4", x"cf", x"e5",
    x"ef", x"10", x"e0", x"22", x"28", x"2e", x"0d", x"fc",
    x"27", x"e6", x"ec", x"2f", x"a4", x"c9", x"11", x"fb",
    x"07", x"f5", x"bc", x"b1", x"bd", x"04", x"02", x"e3",
    x"1c", x"00", x"0a", x"15", x"f9", x"08", x"15", x"0d",
    x"24", x"0b", x"ff", x"11", x"f5", x"19", x"42", x"09",
    x"21", x"16", x"da", x"d8", x"ec", x"c8", x"c7", x"01",
    x"8c", x"a8", x"e1", x"01", x"2a", x"f6", x"9e", x"ed",
    x"df", x"d9", x"e8", x"ec", x"01", x"02", x"07", x"12",
    x"09", x"0a", x"09", x"10", x"0a", x"e8", x"d0", x"d4",
    x"f8", x"ec", x"cb", x"07", x"f8", x"b2", x"e8", x"0e",
    x"10", x"3e", x"3c", x"21", x"de", x"f1", x"1c", x"eb",
    x"f8", x"fe", x"1b", x"fc", x"f4", x"10", x"f3", x"1c",
    x"01", x"fb", x"fc", x"fe", x"06", x"fe", x"fc", x"02",
    x"06", x"fa", x"29", x"38", x"ab", x"98", x"a9", x"dd",
    x"e0", x"c3", x"0e", x"29", x"20", x"e3", x"e4", x"13",
    x"ea", x"05", x"06", x"16", x"f4", x"ff", x"06", x"0f",
    x"0c", x"20", x"e4", x"e5", x"e5", x"f4", x"ef", x"c0",
    x"c0", x"d5", x"09", x"21", x"01", x"2b", x"13", x"25",
    x"ff", x"03", x"1b", x"32", x"3b", x"22", x"ee", x"e8",
    x"24", x"b7", x"d9", x"ea", x"01", x"fd", x"02", x"f1",
    x"de", x"dc", x"18", x"d8", x"fa", x"35", x"ef", x"f5",
    x"00", x"07", x"fc", x"04", x"fd", x"ff", x"09", x"04",
    x"00", x"03", x"02", x"00", x"07", x"08", x"09", x"fc",
    x"02", x"00", x"81", x"e4", x"f2", x"79", x"3d", x"3d",
    x"ff", x"de", x"12", x"cb", x"d5", x"d9", x"e2", x"e1",
    x"e9", x"1c", x"0c", x"d5", x"ec", x"f3", x"f7", x"77",
    x"cc", x"e9", x"11", x"fd", x"da", x"b9", x"cf", x"15",
    x"06", x"b8", x"c7", x"27", x"c6", x"ed", x"be", x"fe",
    x"06", x"bc", x"e9", x"da", x"3a", x"1b", x"fb", x"24",
    x"2b", x"26", x"38", x"e7", x"ea", x"08", x"24", x"ff",
    x"ed", x"22", x"1d", x"cf", x"1d", x"1e", x"ee", x"2b",
    x"26", x"01", x"fc", x"f6", x"1f", x"16", x"0c", x"ff",
    x"10", x"ee", x"06", x"3b", x"0d", x"29", x"ed", x"02",
    x"12", x"c6", x"d7", x"a5", x"ff", x"17", x"f5", x"ad",
    x"cf", x"ee", x"cd", x"df", x"f5", x"e9", x"f2", x"53",
    x"57", x"3d", x"28", x"0e", x"fa", x"11", x"f8", x"11",
    x"91", x"13", x"3d", x"e3", x"00", x"2c", x"ee", x"ce",
    x"f0", x"2f", x"06", x"1b", x"29", x"06", x"f5", x"17",
    x"0b", x"21", x"f7", x"19", x"1c", x"27", x"0a", x"21",
    x"cf", x"d2", x"0d", x"f2", x"ca", x"eb", x"fe", x"e1",
    x"b4", x"36", x"fa", x"12", x"85", x"2a", x"40", x"52",
    x"3f", x"56", x"1c", x"08", x"14", x"e6", x"04", x"1a",
    x"c9", x"ed", x"f2", x"fe", x"dd", x"cc", x"da", x"f1",
    x"27", x"f0", x"d5", x"14", x"eb", x"01", x"1e", x"08",
    x"08", x"e9", x"29", x"fc", x"0c", x"0d", x"10", x"f8",
    x"fa", x"fb", x"cc", x"2e", x"ee", x"b2", x"42", x"f5",
    x"09", x"fe", x"f1", x"01", x"ca", x"ec", x"0a", x"da",
    x"50", x"52", x"59", x"4d", x"39", x"44", x"2c", x"1a",
    x"cc", x"09", x"3f", x"11", x"0b", x"05", x"e2", x"e1",
    x"a9", x"d0", x"dd", x"ce", x"dd", x"0f", x"f4", x"f5",
    x"12", x"26", x"da", x"1c", x"07", x"82", x"e5", x"e0",
    x"1b", x"1b", x"d5", x"c0", x"0e", x"fa", x"aa", x"05",
    x"f7", x"58", x"e5", x"04", x"d0", x"08", x"20", x"0f",
    x"18", x"d5", x"82", x"1f", x"00", x"f0", x"03", x"47",
    x"f0", x"f8", x"42", x"ff", x"f8", x"f1", x"d0", x"dd",
    x"e5", x"05", x"f4", x"0b", x"1a", x"0f", x"01", x"d6",
    x"28", x"1b", x"fc", x"32", x"36", x"ea", x"0e", x"07",
    x"0b", x"fb", x"0e", x"23", x"1d", x"f6", x"ee", x"22",
    x"f2", x"05", x"fd", x"fd", x"fd", x"02", x"04", x"fb",
    x"03", x"03", x"0e", x"09", x"fd", x"07", x"2e", x"23",
    x"21", x"29", x"1c", x"f8", x"d9", x"cc", x"e5", x"c7",
    x"b4", x"3a", x"2a", x"12", x"22", x"fa", x"01", x"42",
    x"18", x"fc", x"5b", x"1d", x"31", x"f7", x"ec", x"d8",
    x"e7", x"f3", x"f5", x"8e", x"50", x"1a", x"e2", x"cd",
    x"ce", x"0c", x"e9", x"d3", x"15", x"0b", x"f2", x"17",
    x"19", x"3a", x"f5", x"fa", x"35", x"06", x"16", x"f6",
    x"ed", x"04", x"09", x"99", x"f8", x"0c", x"07", x"a2",
    x"db", x"f7", x"0d", x"0a", x"17", x"ff", x"e0", x"4a",
    x"f4", x"01", x"f1", x"f8", x"f3", x"d1", x"e2", x"de",
    x"49", x"17", x"21", x"05", x"0a", x"02", x"03", x"0f",
    x"00", x"11", x"0c", x"00", x"24", x"1e", x"33", x"38",
    x"40", x"38", x"03", x"35", x"59", x"26", x"d6", x"08",
    x"da", x"aa", x"d8", x"c4", x"e0", x"f6", x"03", x"09",
    x"06", x"ba", x"29", x"13", x"0e", x"0b", x"07", x"47",
    x"60", x"6c", x"44", x"6a", x"6e", x"82", x"92", x"99",
    x"fd", x"de", x"2f", x"cd", x"c3", x"ea", x"cb", x"ff",
    x"02", x"e8", x"03", x"0e", x"26", x"0b", x"e4", x"fe",
    x"f0", x"e8", x"3b", x"34", x"1a", x"03", x"13", x"1d",
    x"18", x"16", x"34", x"b7", x"1c", x"12", x"ea", x"19",
    x"19", x"23", x"47", x"27", x"07", x"0c", x"0e", x"02",
    x"07", x"11", x"02", x"1b", x"13", x"42", x"09", x"31",
    x"1b", x"01", x"12", x"30", x"04", x"1e", x"1b", x"aa",
    x"fa", x"b2", x"df", x"0b", x"ef", x"e3", x"03", x"ff",
    x"dc", x"1b", x"db", x"cf", x"e6", x"f5", x"f2", x"f6",
    x"fd", x"fe", x"fe", x"ff", x"ff", x"fd", x"04", x"fb",
    x"fd", x"2f", x"15", x"fc", x"08", x"fa", x"ec", x"02",
    x"15", x"f8", x"15", x"45", x"45", x"3a", x"62", x"79",
    x"07", x"34", x"3d", x"13", x"03", x"16", x"e6", x"0b",
    x"01", x"16", x"dc", x"d0", x"34", x"34", x"24", x"da",
    x"e8", x"ec", x"de", x"eb", x"1e", x"41", x"2a", x"44",
    x"47", x"2b", x"fc", x"1c", x"04", x"e2", x"3e", x"03",
    x"e1", x"e8", x"12", x"15", x"f7", x"f6", x"ea", x"24",
    x"0d", x"a2", x"c6", x"b8", x"e7", x"cb", x"f5", x"d8",
    x"05", x"fa", x"04", x"00", x"00", x"fe", x"02", x"0b",
    x"00", x"fc", x"01", x"fb", x"03", x"03", x"02", x"ff",
    x"f9", x"fa", x"c7", x"df", x"ee", x"e9", x"ee", x"cf",
    x"f3", x"ec", x"f8", x"ed", x"cd", x"05", x"e7", x"e1",
    x"eb", x"e9", x"fc", x"00", x"ee", x"e4", x"c5", x"dd",
    x"b3", x"b6", x"03", x"ec", x"eb", x"19", x"09", x"29",
    x"fb", x"38", x"fd", x"1c", x"61", x"f9", x"e5", x"fa",
    x"ff", x"c4", x"ec", x"f5", x"1f", x"1c", x"02", x"4b",
    x"fe", x"f6", x"53", x"17", x"16", x"25", x"e4", x"07",
    x"fd", x"e9", x"11", x"ed", x"df", x"07", x"4e", x"08",
    x"36", x"27", x"1f", x"14", x"0e", x"0e", x"f3", x"ce",
    x"ec", x"c5", x"18", x"f7", x"fa", x"01", x"00", x"e6",
    x"ef", x"03", x"f9", x"f5", x"e2", x"f8", x"14", x"00",
    x"07", x"fe", x"1e", x"f9", x"35", x"1d", x"11", x"76",
    x"2d", x"59", x"4b", x"0c", x"f9", x"06", x"18", x"19",
    x"f6", x"0e", x"22", x"35", x"1c", x"23", x"e3", x"f3",
    x"1e", x"f7", x"1a", x"f8", x"64", x"f2", x"d0", x"39",
    x"0a", x"04", x"fe", x"08", x"f7", x"2a", x"fe", x"1d",
    x"bb", x"da", x"f0", x"f8", x"05", x"21", x"0e", x"21",
    x"24", x"23", x"b7", x"cc", x"09", x"eb", x"08", x"d5",
    x"e5", x"d8", x"1d", x"29", x"0f", x"f0", x"e4", x"e4",
    x"ed", x"02", x"17", x"fb", x"07", x"fc", x"f4", x"e7",
    x"06", x"dd", x"ca", x"f9", x"05", x"e8", x"0b", x"43",
    x"19", x"36", x"ee", x"f8", x"f3", x"ba", x"b0", x"0c",
    x"b8", x"07", x"34", x"18", x"f6", x"f5", x"f1", x"ce",
    x"ea", x"b6", x"eb", x"ff", x"1d", x"22", x"0d", x"e7",
    x"e1", x"f2", x"45", x"0d", x"18", x"2a", x"24", x"ee",
    x"e4", x"ed", x"20", x"24", x"05", x"12", x"0d", x"02",
    x"00", x"0e", x"eb", x"21", x"fe", x"d2", x"ea", x"c5",
    x"fa", x"19", x"e1", x"05", x"0e", x"e0", x"1a", x"2c",
    x"f7", x"38", x"48", x"c2", x"c3", x"c4", x"ec", x"da",
    x"f5", x"14", x"25", x"1f", x"01", x"ce", x"f3", x"05",
    x"f5", x"1f", x"0f", x"05", x"fd", x"8d", x"e6", x"e8",
    x"cd", x"d7", x"ec", x"fd", x"fe", x"31", x"f5", x"f8",
    x"43", x"ff", x"17", x"06", x"2b", x"1c", x"1d", x"18",
    x"fe", x"c0", x"f3", x"e1", x"15", x"e7", x"4a", x"35",
    x"00", x"b7", x"dc", x"16", x"1a", x"3b", x"1c", x"1c",
    x"11", x"fe", x"fb", x"fb", x"fb", x"03", x"00", x"00",
    x"fe", x"03", x"fd", x"13", x"e4", x"d2", x"ec", x"b5",
    x"10", x"02", x"13", x"ff", x"d9", x"0a", x"e5", x"e9",
    x"e6", x"d7", x"ea", x"c3", x"7c", x"9c", x"be", x"d1",
    x"b6", x"f8", x"ea", x"df", x"ad", x"e8", x"d5", x"f8",
    x"07", x"02", x"17", x"05", x"d9", x"ce", x"d1", x"be",
    x"c0", x"ff", x"07", x"fb", x"31", x"18", x"cf", x"ee",
    x"c5", x"91", x"09", x"02", x"2f", x"d7", x"06", x"ff",
    x"04", x"c9", x"80", x"f2", x"da", x"ce", x"f2", x"2c",
    x"18", x"ec", x"10", x"0d", x"fd", x"ee", x"17", x"ab",
    x"1b", x"19", x"f5", x"03", x"0f", x"01", x"14", x"02",
    x"b4", x"be", x"ad", x"fb", x"fe", x"ff", x"fc", x"fb",
    x"fb", x"01", x"fb", x"01", x"14", x"04", x"17", x"35",
    x"f7", x"20", x"07", x"0e", x"39", x"f8", x"c5", x"c3",
    x"32", x"16", x"f5", x"24", x"ed", x"35", x"07", x"de",
    x"b9", x"ed", x"fa", x"fb", x"1e", x"18", x"2e", x"e5",
    x"e9", x"21", x"19", x"0c", x"05", x"11", x"26", x"0f",
    x"c6", x"c0", x"a2", x"cc", x"d3", x"f7", x"e8", x"ea",
    x"f7", x"1a", x"03", x"0d", x"a7", x"b5", x"f3", x"d3",
    x"c6", x"32", x"e0", x"f9", x"dc", x"f3", x"f7", x"f2",
    x"ef", x"19", x"2e", x"07", x"f3", x"83", x"e2", x"fd",
    x"e7", x"10", x"05", x"f1", x"0e", x"11", x"06", x"08",
    x"0a", x"02", x"0d", x"0c", x"04", x"e5", x"ec", x"f7",
    x"e4", x"d9", x"19", x"22", x"f5", x"00", x"fa", x"f7",
    x"e0", x"c2", x"34", x"1a", x"f0", x"24", x"05", x"e3",
    x"cf", x"f5", x"bb", x"ef", x"00", x"15", x"35", x"20",
    x"fb", x"fb", x"fc", x"02", x"06", x"00", x"fd", x"fe",
    x"03", x"d3", x"d9", x"d4", x"fc", x"0d", x"f0", x"02",
    x"00", x"01", x"f7", x"0e", x"17", x"06", x"1c", x"1c",
    x"47", x"25", x"0a", x"d0", x"e3", x"ed", x"e3", x"f8",
    x"f5", x"f5", x"dc", x"fb", x"35", x"21", x"d2", x"fc",
    x"0e", x"1c", x"ea", x"a2", x"f0", x"dc", x"bf", x"06",
    x"fe", x"df", x"01", x"12", x"0b", x"f7", x"3a", x"25",
    x"c9", x"d1", x"b9", x"eb", x"dc", x"d7", x"14", x"db",
    x"00", x"ca", x"c4", x"da", x"f5", x"a9", x"cf", x"f9",
    x"04", x"03", x"00", x"ff", x"03", x"04", x"00", x"05",
    x"01", x"00", x"00", x"ff", x"00", x"02", x"fa", x"02",
    x"fc", x"ff", x"06", x"e7", x"4d", x"34", x"f8", x"11",
    x"f1", x"f7", x"f6", x"c3", x"07", x"f3", x"be", x"b9",
    x"fa", x"0a", x"06", x"fb", x"b9", x"df", x"dc", x"ce",
    x"cc", x"e8", x"de", x"f1", x"15", x"fa", x"c6", x"f9",
    x"11", x"11", x"17", x"06", x"ef", x"e2", x"1e", x"f9",
    x"f6", x"10", x"d9", x"09", x"c2", x"ba", x"c9", x"e0",
    x"a7", x"56", x"00", x"f9", x"d2", x"4d", x"2b", x"fd",
    x"d7", x"d4", x"fb", x"08", x"e4", x"f9", x"3c", x"cd",
    x"1d", x"b4", x"dc", x"05", x"e9", x"d6", x"fb", x"e7",
    x"df", x"cc", x"b8", x"cf", x"af", x"d9", x"e5", x"fb",
    x"27", x"08", x"17", x"45", x"23", x"40", x"23", x"01",
    x"0b", x"fe", x"0b", x"0f", x"01", x"e5", x"e2", x"e2",
    x"23", x"16", x"10", x"ea", x"18", x"d5", x"ba", x"e0",
    x"fb", x"31", x"22", x"13", x"07", x"12", x"ea", x"cf",
    x"da", x"12", x"0c", x"ff", x"3d", x"20", x"f6", x"df",
    x"f2", x"08", x"d5", x"f4", x"f6", x"f0", x"fc", x"08",
    x"0c", x"dd", x"e4", x"3b", x"0a", x"d9", x"03", x"fc",
    x"10", x"e9", x"04", x"0c", x"15", x"13", x"dd", x"e9",
    x"0f", x"dc", x"cf", x"d5", x"e7", x"9a", x"bf", x"f4",
    x"e9", x"e1", x"d4", x"ec", x"13", x"04", x"ca", x"05",
    x"fa", x"e7", x"f1", x"08", x"fb", x"f5", x"ff", x"f1",
    x"15", x"e2", x"de", x"fb", x"fa", x"0e", x"18", x"fa",
    x"f3", x"0c", x"f9", x"f2", x"f3", x"e9", x"03", x"fe",
    x"e8", x"1d", x"e3", x"11", x"f2", x"0c", x"fd", x"fe",
    x"1f", x"05", x"17", x"e9", x"06", x"10", x"08", x"e7",
    x"02", x"f3", x"1b", x"0c", x"f7", x"bc", x"20", x"ed",
    x"e4", x"c9", x"13", x"f5", x"1d", x"0e", x"1f", x"20",
    x"16", x"08", x"01", x"cc", x"e9", x"17", x"f2", x"04",
    x"f8", x"e3", x"f0", x"01", x"d6", x"e9", x"eb", x"f4",
    x"da", x"03", x"02", x"f6", x"1d", x"0f", x"ce", x"0d",
    x"0c", x"cd", x"05", x"e5", x"f5", x"ec", x"e9", x"06",
    x"e0", x"f4", x"fb", x"e1", x"03", x"01", x"f9", x"ff",
    x"0d", x"0f", x"e9", x"23", x"f8", x"ec", x"0f", x"f4",
    x"b9", x"de", x"ec", x"da", x"f6", x"da", x"10", x"16",
    x"2a", x"36", x"d4", x"03", x"3a", x"e3", x"20", x"28",
    x"11", x"03", x"fd", x"fe", x"fe", x"05", x"fb", x"06",
    x"fe", x"01", x"f9", x"d4", x"0e", x"ec", x"e4", x"13",
    x"13", x"e8", x"f4", x"0a", x"fe", x"19", x"0a", x"13",
    x"09", x"1e", x"01", x"0d", x"0f", x"e3", x"29", x"03",
    x"0e", x"34", x"02", x"22", x"29", x"1f", x"02", x"e7",
    x"12", x"07", x"f3", x"ed", x"22", x"ea", x"32", x"ee",
    x"ec", x"28", x"28", x"e2", x"01", x"fd", x"13", x"19",
    x"0f", x"fb", x"0e", x"fd", x"0e", x"fa", x"fd", x"ed",
    x"36", x"ec", x"d4", x"3f", x"13", x"e0", x"f7", x"ec",
    x"ed", x"fb", x"c1", x"1c", x"0e", x"1c", x"1c", x"09",
    x"fc", x"1a", x"fc", x"05", x"e8", x"21", x"2c", x"0b",
    x"d5", x"05", x"e5", x"02", x"00", x"fc", x"01", x"05",
    x"03", x"00", x"03", x"04", x"24", x"11", x"11", x"0c",
    x"ff", x"04", x"03", x"f8", x"e2", x"1f", x"17", x"28",
    x"0d", x"e2", x"f1", x"01", x"0d", x"3b", x"0b", x"dc",
    x"d8", x"f1", x"2a", x"ee", x"0d", x"0f", x"02", x"04",
    x"e0", x"30", x"f9", x"f8", x"ff", x"fa", x"fd", x"0e",
    x"04", x"ba", x"18", x"1c", x"cd", x"c5", x"11", x"cd",
    x"c3", x"03", x"cf", x"de", x"0b", x"07", x"1a", x"12",
    x"f5", x"00", x"ec", x"f7", x"ee", x"e0", x"cb", x"f2",
    x"17", x"da", x"b9", x"16", x"0e", x"e0", x"36", x"0d",
    x"04", x"0e", x"08", x"09", x"00", x"f4", x"f5", x"00",
    x"04", x"03", x"01", x"03", x"fb", x"00", x"07", x"06",
    x"00", x"fe", x"d8", x"ec", x"2d", x"ec", x"43", x"cb",
    x"ec", x"0e", x"d1", x"fc", x"ee", x"d0", x"f2", x"1f",
    x"fb", x"16", x"f8", x"15", x"ec", x"1b", x"f3", x"fe",
    x"05", x"ff", x"fb", x"00", x"01", x"01", x"03", x"02",
    x"01", x"e0", x"bc", x"da", x"e2", x"e4", x"f3", x"2a",
    x"1a", x"13", x"ed", x"ec", x"10", x"06", x"1d", x"0c",
    x"fb", x"25", x"1b", x"f3", x"ce", x"d6", x"f8", x"0a",
    x"e5", x"24", x"02", x"ec", x"f0", x"06", x"12", x"03",
    x"14", x"1d", x"d6", x"14", x"02", x"f4", x"17", x"27",
    x"fe", x"f0", x"d9", x"06", x"06", x"07", x"09", x"33",
    x"0b", x"2a", x"fd", x"19", x"0f", x"fc", x"0f", x"f2",
    x"1c", x"ff", x"ff", x"e0", x"0a", x"13", x"ee", x"09",
    x"fb", x"04", x"04", x"fc", x"fd", x"05", x"01", x"fb",
    x"fd", x"00", x"00", x"fc", x"03", x"03", x"ff", x"01",
    x"ff", x"03", x"35", x"08", x"15", x"0a", x"14", x"dd",
    x"22", x"fc", x"f1", x"18", x"db", x"e1", x"2f", x"ea",
    x"cc", x"08", x"f2", x"da", x"05", x"06", x"0b", x"e7",
    x"ef", x"31", x"04", x"00", x"ea", x"df", x"e5", x"f8",
    x"e4", x"e8", x"ed", x"05", x"0a", x"ed", x"11", x"1f",
    x"cd", x"27", x"13", x"03", x"05", x"c9", x"dc", x"06",
    x"14", x"e1", x"ed", x"0d", x"cc", x"03", x"d0", x"22",
    x"0b", x"04", x"c0", x"0f", x"d7", x"cb", x"1b", x"fa",
    x"04", x"d7", x"fb", x"31", x"c0", x"fc", x"f7", x"07",
    x"04", x"de", x"0f", x"ec", x"cb", x"0b", x"e3", x"dd",
    x"ff", x"f8", x"e4", x"f7", x"ea", x"e8", x"f6", x"0e",
    x"03", x"f8", x"eb", x"cc", x"e4", x"03", x"17", x"36",
    x"00", x"15", x"0a", x"18", x"02", x"26", x"3e", x"23",
    x"10", x"0a", x"f5", x"18", x"17", x"f1", x"1d", x"0d",
    x"08", x"28", x"07", x"fc", x"1c", x"eb", x"ce", x"3a",
    x"10", x"2b", x"0c", x"06", x"e9", x"02", x"f2", x"06",
    x"b5", x"b3", x"f3", x"e2", x"fe", x"2d", x"0c", x"25",
    x"40", x"47", x"f0", x"f3", x"72", x"df", x"08", x"64",
    x"0f", x"10", x"2f", x"37", x"2c", x"11", x"3a", x"3e",
    x"0b", x"26", x"15", x"d2", x"e3", x"f8", x"35", x"1a",
    x"fa", x"92", x"84", x"b0", x"d5", x"19", x"36", x"0c",
    x"3b", x"4f", x"18", x"1f", x"19", x"2a", x"36", x"ef",
    x"ff", x"ea", x"2f", x"e5", x"f3", x"04", x"2b", x"e2",
    x"dc", x"b3", x"ac", x"cd", x"eb", x"91", x"ae", x"f9",
    x"02", x"21", x"8a", x"9d", x"45", x"fb", x"e2", x"e1",
    x"14", x"35", x"0f", x"f5", x"13", x"0b", x"f2", x"ff",
    x"17", x"42", x"39", x"1b", x"e2", x"ea", x"10", x"4d",
    x"0d", x"12", x"54", x"0e", x"ff", x"2e", x"bc", x"d6",
    x"46", x"38", x"f4", x"e0", x"d1", x"c7", x"31", x"d1",
    x"c7", x"33", x"db", x"cd", x"74", x"e5", x"25", x"bd",
    x"29", x"22", x"38", x"24", x"3a", x"30", x"2c", x"02",
    x"31", x"14", x"0e", x"fe", x"e9", x"fc", x"14", x"02",
    x"e7", x"fa", x"e6", x"d8", x"bc", x"db", x"ff", x"81",
    x"f6", x"14", x"74", x"4f", x"0a", x"0f", x"02", x"d8",
    x"b5", x"df", x"dc", x"b7", x"e3", x"e3", x"f0", x"fc",
    x"50", x"fd", x"fb", x"01", x"fd", x"02", x"fd", x"fe",
    x"01", x"01", x"53", x"77", x"5c", x"1b", x"e8", x"ca",
    x"ee", x"ef", x"06", x"0d", x"f2", x"ef", x"27", x"f2",
    x"e7", x"11", x"f3", x"fd", x"3c", x"fb", x"0e", x"1a",
    x"26", x"01", x"02", x"0f", x"f5", x"05", x"ff", x"fe",
    x"10", x"fd", x"eb", x"23", x"11", x"fc", x"e1", x"21",
    x"06", x"a3", x"c4", x"f7", x"29", x"14", x"41", x"01",
    x"e9", x"fe", x"14", x"0f", x"1e", x"45", x"39", x"2f",
    x"27", x"e0", x"f9", x"d9", x"06", x"19", x"ec", x"43",
    x"28", x"fc", x"01", x"14", x"c1", x"dc", x"18", x"d8",
    x"f2", x"f7", x"24", x"13", x"20", x"33", x"ee", x"f1",
    x"0d", x"de", x"e4", x"0a", x"06", x"07", x"0b", x"08",
    x"ff", x"0f", x"07", x"03", x"12", x"ff", x"3f", x"da",
    x"0f", x"0e", x"d2", x"ec", x"24", x"e5", x"fe", x"c0",
    x"80", x"92", x"b1", x"1c", x"db", x"ce", x"1e", x"1f",
    x"37", x"e6", x"fd", x"17", x"d9", x"ee", x"21", x"d4",
    x"ff", x"07", x"cc", x"fc", x"07", x"11", x"fb", x"d3",
    x"1c", x"2c", x"18", x"c4", x"e6", x"07", x"f7", x"fc",
    x"26", x"4d", x"03", x"f9", x"16", x"28", x"18", x"04",
    x"de", x"00", x"e3", x"11", x"ff", x"ad", x"ae", x"cf",
    x"a4", x"d2", x"ce", x"f0", x"fd", x"16", x"ef", x"00",
    x"f5", x"3b", x"f5", x"f8", x"fa", x"03", x"05", x"ff",
    x"00", x"fa", x"fb", x"f5", x"fd", x"35", x"1d", x"31",
    x"0c", x"b9", x"b0", x"dd", x"c9", x"e1", x"46", x"03",
    x"f3", x"f4", x"39", x"28", x"74", x"37", x"21", x"62",
    x"0c", x"e1", x"0c", x"ec", x"e5", x"31", x"fc", x"0b",
    x"05", x"fe", x"03", x"fb", x"06", x"fd", x"ff", x"fd",
    x"01", x"fd", x"1a", x"1a", x"23", x"0d", x"30", x"08",
    x"b6", x"d4", x"fd", x"9f", x"c4", x"c1", x"06", x"eb",
    x"0f", x"fe", x"ee", x"5c", x"eb", x"e8", x"01", x"ee",
    x"0f", x"15", x"f2", x"16", x"71", x"67", x"56", x"ee",
    x"e0", x"e1", x"e2", x"f5", x"f3", x"83", x"dd", x"f4",
    x"f9", x"25", x"20", x"2c", x"1e", x"30", x"33", x"f8",
    x"04", x"39", x"f7", x"d8", x"03", x"f1", x"1a", x"56",
    x"2f", x"2f", x"21", x"20", x"31", x"ee", x"25", x"1b",
    x"02", x"fe", x"fa", x"fe", x"03", x"03", x"fd", x"fc",
    x"06", x"04", x"06", x"06", x"fc", x"01", x"fd", x"fc",
    x"ff", x"01", x"ee", x"c0", x"f7", x"fb", x"0c", x"f4",
    x"52", x"03", x"fe", x"f4", x"fc", x"f6", x"02", x"f1",
    x"ec", x"ff", x"ff", x"05", x"3f", x"3f", x"39", x"31",
    x"3e", x"01", x"bb", x"ee", x"26", x"06", x"06", x"2f",
    x"f5", x"fd", x"09", x"5b", x"3d", x"e3", x"4a", x"e3",
    x"18", x"f7", x"cd", x"25", x"ed", x"da", x"0f", x"fb",
    x"d5", x"e0", x"e9", x"a9", x"cd", x"02", x"99", x"ab",
    x"cf", x"96", x"ed", x"a6", x"60", x"de", x"15", x"f9",
    x"09", x"07", x"39", x"42", x"11", x"28", x"27", x"10",
    x"26", x"17", x"f2", x"0f", x"3c", x"13", x"39", x"43",
    x"33", x"f2", x"ff", x"33", x"1a", x"0a", x"01", x"1e",
    x"2e", x"df", x"fc", x"02", x"3c", x"ff", x"ae", x"f6",
    x"05", x"02", x"4f", x"25", x"1e", x"17", x"f4", x"ed",
    x"0c", x"b3", x"10", x"65", x"f7", x"06", x"d3", x"0e",
    x"0b", x"88", x"16", x"16", x"07", x"f5", x"16", x"eb",
    x"08", x"e5", x"96", x"ce", x"ce", x"e2", x"0a", x"0b",
    x"f8", x"f7", x"01", x"ff", x"e5", x"13", x"03", x"de",
    x"22", x"c8", x"d1", x"d4", x"e4", x"cf", x"e0", x"c2",
    x"d8", x"d4", x"f7", x"0d", x"2e", x"12", x"f4", x"18",
    x"02", x"f0", x"37", x"ef", x"e6", x"e3", x"0b", x"db",
    x"f9", x"1f", x"1a", x"03", x"fd", x"2c", x"d9", x"09",
    x"16", x"cd", x"b6", x"d5", x"c2", x"1c", x"0e", x"b3",
    x"15", x"07", x"18", x"ff", x"16", x"30", x"1d", x"20",
    x"06", x"fe", x"11", x"1a", x"0b", x"3c", x"31", x"1d",
    x"18", x"2d", x"f1", x"e4", x"bf", x"18", x"c4", x"b2",
    x"f5", x"d0", x"bb", x"10", x"b7", x"70", x"f2", x"b3",
    x"a1", x"2e", x"ef", x"eb", x"16", x"f2", x"0f", x"0d",
    x"1e", x"e1", x"0a", x"ec", x"f7", x"3d", x"d9", x"04",
    x"00", x"00", x"f3", x"3b", x"0f", x"19", x"05", x"17",
    x"1b", x"fb", x"2d", x"31", x"5d", x"da", x"f1", x"1e",
    x"d7", x"00", x"06", x"f2", x"07", x"0d", x"e7", x"6d",
    x"04", x"00", x"ab", x"28", x"16", x"ee", x"22", x"12",
    x"28", x"20", x"40", x"45", x"47", x"49", x"49", x"f1",
    x"05", x"2d", x"eb", x"ed", x"c4", x"ea", x"e3", x"de",
    x"0e", x"fd", x"d3", x"01", x"dc", x"ce", x"fb", x"e6",
    x"e3", x"00", x"fd", x"fe", x"fd", x"03", x"fc", x"03",
    x"fc", x"01", x"1a", x"0d", x"10", x"1f", x"09", x"ef",
    x"11", x"f3", x"0f", x"f5", x"e1", x"0b", x"ee", x"0e",
    x"2d", x"1f", x"f2", x"f2", x"13", x"b8", x"b0", x"0a",
    x"eb", x"9a", x"f2", x"e7", x"aa", x"13", x"f6", x"11",
    x"f7", x"eb", x"ed", x"c1", x"f0", x"fc", x"0a", x"13",
    x"33", x"36", x"fb", x"1d", x"cd", x"d3", x"e5", x"00",
    x"d3", x"e3", x"cc", x"07", x"f1", x"c5", x"db", x"bb",
    x"e2", x"a9", x"04", x"2c", x"c8", x"07", x"18", x"2a",
    x"24", x"e0", x"ad", x"aa", x"f5", x"e0", x"d6", x"fa",
    x"08", x"08", x"f2", x"18", x"eb", x"ec", x"02", x"d3",
    x"f7", x"1c", x"f5", x"fc", x"f9", x"fe", x"fe", x"09",
    x"0e", x"03", x"ff", x"02", x"16", x"39", x"44", x"f4",
    x"05", x"1b", x"d2", x"03", x"cd", x"0d", x"20", x"3a",
    x"f3", x"08", x"09", x"e3", x"ee", x"c9", x"23", x"f6",
    x"11", x"0a", x"f0", x"0f", x"1c", x"0d", x"fe", x"2e",
    x"fa", x"e6", x"f7", x"fa", x"d8", x"01", x"f7", x"a9",
    x"0e", x"38", x"2c", x"0e", x"21", x"46", x"34", x"49",
    x"58", x"15", x"f8", x"e6", x"f0", x"1f", x"bd", x"09",
    x"3d", x"db", x"1f", x"f4", x"05", x"22", x"23", x"3c",
    x"27", x"17", x"2f", x"e1", x"e2", x"ca", x"06", x"98",
    x"99", x"bf", x"6a", x"62", x"08", x"0a", x"14", x"0d",
    x"08", x"02", x"01", x"01", x"fa", x"f5", x"c2", x"d4",
    x"ec", x"d3", x"be", x"f2", x"d3", x"af", x"f8", x"0e",
    x"1d", x"15", x"24", x"27", x"04", x"34", x"30", x"cf",
    x"0f", x"18", x"f8", x"47", x"45", x"41", x"45", x"33",
    x"00", x"05", x"ff", x"ff", x"00", x"04", x"05", x"01",
    x"05", x"0b", x"ea", x"e1", x"f8", x"d5", x"d8", x"d3",
    x"db", x"f0", x"d4", x"d1", x"c3", x"b2", x"da", x"bf",
    x"be", x"f5", x"a1", x"14", x"db", x"e0", x"01", x"ce",
    x"d7", x"e1", x"b4", x"bb", x"f5", x"de", x"85", x"ff",
    x"f3", x"d6", x"06", x"fb", x"e6", x"bd", x"b8", x"dd",
    x"e6", x"be", x"cd", x"f2", x"df", x"d5", x"e8", x"ef",
    x"38", x"00", x"dd", x"c8", x"07", x"d4", x"ef", x"20",
    x"09", x"1e", x"19", x"10", x"32", x"06", x"2d", x"4d",
    x"fd", x"fe", x"06", x"fb", x"03", x"03", x"ff", x"06",
    x"fc", x"fb", x"03", x"ff", x"fd", x"04", x"03", x"01",
    x"fc", x"fe", x"12", x"03", x"02", x"01", x"04", x"01",
    x"1e", x"1c", x"08", x"2e", x"0d", x"29", x"13", x"20",
    x"4c", x"23", x"3e", x"59", x"14", x"29", x"20", x"0b",
    x"1b", x"1c", x"0a", x"1c", x"f4", x"24", x"41", x"2a",
    x"2b", x"38", x"05", x"d7", x"f2", x"fd", x"36", x"38",
    x"22", x"3c", x"39", x"41", x"0f", x"1e", x"30", x"ee",
    x"f8", x"1b", x"39", x"d8", x"12", x"5c", x"32", x"fd",
    x"13", x"ff", x"2a", x"00", x"e7", x"01", x"2f", x"07",
    x"fe", x"e6", x"0e", x"25", x"c1", x"df", x"f5", x"03",
    x"f5", x"0f", x"e4", x"0f", x"22", x"f4", x"02", x"22",
    x"fd", x"f8", x"12", x"1e", x"14", x"08", x"18", x"04",
    x"11", x"32", x"2a", x"2a", x"12", x"0b", x"a4", x"01",
    x"e5", x"c1", x"dc", x"c1", x"10", x"e2", x"15", x"0d",
    x"1c", x"07", x"fc", x"cb", x"a4", x"90", x"17", x"37",
    x"1c", x"1c", x"dc", x"ef", x"10", x"c9", x"ef", x"08",
    x"11", x"11", x"1b", x"10", x"22", x"24", x"19", x"33",
    x"fd", x"fd", x"fb", x"ff", x"04", x"01", x"fa", x"fc",
    x"ff", x"fc", x"fa", x"fe", x"f7", x"fe", x"fe", x"00",
    x"fe", x"01", x"fc", x"fb", x"02", x"fa", x"00", x"02",
    x"ff", x"fd", x"03", x"00", x"f9", x"f9", x"fb", x"02",
    x"f9", x"fa", x"fc", x"f9", x"05", x"fb", x"00", x"fa",
    x"ff", x"fd", x"ff", x"fa", x"ff", x"fa", x"fb", x"fb",
    x"fd", x"ff", x"01", x"02", x"ff", x"03", x"fb", x"fe",
    x"00", x"00", x"fe", x"f9", x"fa", x"fc", x"fc", x"04",
    x"fc", x"00", x"f7", x"04", x"01", x"01", x"01", x"fa",
    x"fa", x"02", x"02", x"fe", x"fc", x"02", x"03", x"fd",
    x"fa", x"fb", x"f9", x"05", x"00", x"fb", x"01", x"fe",
    x"02", x"fb", x"03", x"01", x"f8", x"fb", x"fb", x"fb",
    x"00", x"ff", x"fa", x"fe", x"fc", x"01", x"fd", x"f8",
    x"f8", x"04", x"fe", x"fa", x"00", x"fe", x"f9", x"00",
    x"fe", x"fe", x"fa", x"fc", x"fe", x"fa", x"fb", x"03",
    x"00", x"ff", x"04", x"fa", x"f8", x"f7", x"02", x"02",
    x"fc", x"fe", x"00", x"fd", x"03", x"fd", x"fb", x"f7",
    x"02", x"01", x"fc", x"ff", x"f9", x"ff", x"01", x"fb",
    x"00", x"03", x"fe", x"04", x"fd", x"00", x"03", x"00",
    x"00", x"04", x"fb", x"fe", x"00", x"fe", x"00", x"fe",
    x"fb", x"fe", x"fc", x"fd", x"00", x"fa", x"fc", x"04",
    x"02", x"fc", x"fa", x"fb", x"fa", x"04", x"00", x"fd",
    x"fb", x"ff", x"03", x"ff", x"f8", x"00", x"02", x"fe",
    x"ff", x"fa", x"fc", x"fe", x"fd", x"00", x"fb", x"fa",
    x"fe", x"fe", x"ff", x"fd", x"02", x"fd", x"04", x"ff",
    x"ff", x"02", x"02", x"ff", x"fe", x"ff", x"04", x"fd",
    x"01", x"00", x"f8", x"fc", x"fc", x"fe", x"fc", x"ff",
    x"05", x"04", x"fc", x"fd", x"06", x"fd", x"04", x"ff",
    x"fd", x"fe", x"f8", x"fe", x"03", x"ff", x"f8", x"00",
    x"ff", x"04", x"fe", x"00", x"00", x"fb", x"fe", x"03",
    x"08", x"02", x"04", x"05", x"fd", x"fe", x"fb", x"00",
    x"00", x"05", x"fc", x"03", x"02", x"fc", x"00", x"f9",
    x"f7", x"fa", x"02", x"fb", x"ff", x"f7", x"02", x"fa",
    x"f8", x"02", x"fc", x"01", x"00", x"fe", x"00", x"fc",
    x"00", x"fb", x"05", x"fd", x"fc", x"fb", x"ff", x"01",
    x"fa", x"02", x"f8", x"f7", x"fd", x"fc", x"fa", x"02",
    x"fb", x"00", x"02", x"fd", x"f9", x"fb", x"fc", x"02",
    x"00", x"fd", x"fd", x"f9", x"00", x"06", x"05", x"02",
    x"00", x"03", x"04", x"fb", x"02", x"fd", x"ff", x"fe",
    x"04", x"fe", x"fc", x"fc", x"00", x"f8", x"00", x"f9",
    x"02", x"01", x"01", x"fe", x"01", x"01", x"00", x"fb",
    x"02", x"ff", x"fe", x"ff", x"02", x"fc", x"00", x"ff",
    x"f7", x"f7", x"01", x"01", x"00", x"01", x"fa", x"01",
    x"fa", x"00", x"fb", x"fc", x"fc", x"fc", x"fa", x"fc",
    x"ff", x"03", x"ff", x"04", x"fa", x"fb", x"04", x"fd",
    x"fe", x"03", x"fc", x"01", x"02", x"fa", x"03", x"04",
    x"00", x"00", x"ff", x"03", x"fd", x"fa", x"fc", x"f9",
    x"fc", x"00", x"fb", x"fc", x"fa", x"ff", x"f8", x"03",
    x"fc", x"01", x"fc", x"03", x"02", x"fa", x"fa", x"00",
    x"00", x"02", x"fe", x"ff", x"02", x"fb", x"01", x"fb",
    x"04", x"03", x"f7", x"f7", x"fd", x"04", x"02", x"ff",
    x"fa", x"fb", x"04", x"01", x"fb", x"fa", x"fc", x"04",
    x"03", x"04", x"03", x"00", x"06", x"fd", x"fc", x"fb",
    x"00", x"fd", x"ff", x"00", x"fa", x"07", x"ff", x"02",
    x"03", x"04", x"fc", x"04", x"04", x"04", x"02", x"02",
    x"fd", x"00", x"ff", x"fd", x"00", x"00", x"00", x"04",
    x"03", x"fd", x"f9", x"04", x"fd", x"fe", x"03", x"fc",
    x"fb", x"01", x"fd", x"fe", x"fa", x"fc", x"f8", x"ff",
    x"fd", x"00", x"ff", x"04", x"fa", x"fb", x"ff", x"ff",
    x"ff", x"ff", x"01", x"fb", x"fb", x"ff", x"fb", x"00",
    x"f8", x"00", x"fe", x"fa", x"fa", x"01", x"00", x"02",
    x"fb", x"fc", x"03", x"03", x"00", x"f9", x"00", x"ff",
    x"02", x"fe", x"fe", x"fb", x"fd", x"fb", x"00", x"01",
    x"f9", x"fc", x"fc", x"03", x"ff", x"fa", x"fd", x"fc",
    x"fc", x"00", x"f9", x"ff", x"f8", x"fb", x"f7", x"00",
    x"ff", x"01", x"f9", x"fe", x"fc", x"00", x"ff", x"02",
    x"fa", x"fa", x"01", x"f8", x"fd", x"fc", x"fa", x"01",
    x"ff", x"04", x"fc", x"fa", x"fd", x"fa", x"01", x"fe",
    x"02", x"fc", x"fd", x"02", x"fd", x"fc", x"fc", x"fa",
    x"f8", x"fb", x"fa", x"fd", x"fa", x"f8", x"04", x"05",
    x"02", x"fc", x"ff", x"06", x"ff", x"fd", x"02", x"fe",
    x"fd", x"02", x"ff", x"f6", x"00", x"f9", x"fd", x"01",
    x"01", x"ff", x"fe", x"fb", x"ff", x"fb", x"00", x"04",
    x"fc", x"f9", x"fe", x"fc", x"03", x"ff", x"fd", x"fc",
    x"02", x"ff", x"00", x"fb", x"00", x"fa", x"fc", x"fb",
    x"fe", x"fb", x"02", x"fb", x"fa", x"fd", x"fd", x"fe",
    x"f7", x"fd", x"fe", x"f9", x"fd", x"ff", x"01", x"fb",
    x"fa", x"04", x"01", x"02", x"02", x"fd", x"04", x"03",
    x"02", x"04", x"fe", x"00", x"02", x"00", x"00", x"04",
    x"fc", x"fe", x"fd", x"fc", x"fc", x"01", x"ff", x"02",
    x"02", x"01", x"fe", x"01", x"fa", x"03", x"01", x"ff",
    x"fd", x"01", x"ff", x"fa", x"fb", x"ff", x"fb", x"fb",
    x"03", x"00", x"fd", x"ff", x"fb", x"ff", x"00", x"fb",
    x"01", x"fb", x"fd", x"03", x"fb", x"fe", x"fb", x"01",
    x"fd", x"01", x"fd", x"01", x"fe", x"02", x"00", x"02",
    x"00", x"01", x"ff", x"f9", x"05", x"fd", x"01", x"03",
    x"02", x"fd", x"03", x"fe", x"ff", x"fc", x"fb", x"fb",
    x"ff", x"02", x"00", x"fb", x"f9", x"f6", x"fd", x"03",
    x"02", x"fb", x"fd", x"03", x"fe", x"fb", x"fa", x"fe",
    x"fb", x"fa", x"fa", x"fb", x"fe", x"fb", x"02", x"fb",
    x"fd", x"fc", x"02", x"fb", x"fe", x"04", x"04", x"00",
    x"fb", x"03", x"fb", x"ff", x"fb", x"01", x"00", x"05",
    x"04", x"fb", x"fc", x"01", x"03", x"fa", x"03", x"fc",
    x"fe", x"01", x"01", x"03", x"02", x"01", x"01", x"01",
    x"f8", x"02", x"fa", x"fc", x"f9", x"fe", x"fc", x"fc",
    x"fc", x"ff", x"01", x"02", x"fc", x"fc", x"fe", x"01",
    x"fd", x"02", x"fe", x"03", x"fc", x"01", x"ff", x"01",
    x"ff", x"00", x"01", x"fe", x"ff", x"fd", x"fe", x"04",
    x"fb", x"02", x"00", x"01", x"fc", x"00", x"02", x"03",
    x"fb", x"01", x"fa", x"fc", x"02", x"01", x"00", x"00",
    x"00", x"fb", x"fa", x"fd", x"fa", x"fb", x"fb", x"02",
    x"00", x"fa", x"02", x"02", x"fb", x"fc", x"ff", x"00",
    x"fc", x"01", x"ff", x"fd", x"00", x"03", x"02", x"fd",
    x"ff", x"fe", x"00", x"01", x"01", x"fe", x"01", x"04",
    x"03", x"ff", x"ff", x"fc", x"fe", x"fb", x"03", x"02",
    x"fa", x"fd", x"04", x"00", x"03", x"fe", x"ff", x"04",
    x"06", x"00", x"03", x"ff", x"02", x"02", x"fb", x"01",
    x"fd", x"00", x"fb", x"fc", x"fb", x"fd", x"fd", x"fc",
    x"ff", x"fb", x"fb", x"00", x"fe", x"fd", x"fa", x"fc",
    x"fe", x"00", x"fa", x"f9", x"fb", x"00", x"00", x"fa",
    x"03", x"00", x"fe", x"03", x"fd", x"fd", x"ff", x"fe",
    x"fe", x"ff", x"fc", x"03", x"fc", x"02", x"f9", x"00",
    x"f9", x"00", x"fc", x"fb", x"02", x"01", x"00", x"03",
    x"04", x"01", x"00", x"03", x"fc", x"00", x"fb", x"fc",
    x"fa", x"02", x"fd", x"00", x"fd", x"fb", x"fc", x"fb",
    x"00", x"fe", x"00", x"00", x"fe", x"02", x"fe", x"f6",
    x"fe", x"fa", x"ff", x"03", x"01", x"f9", x"fa", x"ff",
    x"00", x"fc", x"00", x"03", x"ff", x"fe", x"02", x"00",
    x"00", x"02", x"fd", x"04", x"01", x"02", x"05", x"fb",
    x"fa", x"fc", x"fb", x"00", x"02", x"ff", x"fd", x"ff",
    x"01", x"ff", x"fe", x"01", x"fb", x"fe", x"fd", x"fc",
    x"fe", x"04", x"01", x"00", x"03", x"fd", x"04", x"01",
    x"fb", x"fc", x"00", x"fb", x"f8", x"fd", x"05", x"fd",
    x"00", x"ff", x"00", x"00", x"ff", x"fa", x"fd", x"02",
    x"fd", x"01", x"ff", x"00", x"fe", x"fa", x"fa", x"04",
    x"fe", x"04", x"02", x"01", x"ff", x"00", x"00", x"fe",
    x"ff", x"fc", x"ff", x"fb", x"03", x"03", x"ff", x"fd",
    x"05", x"01", x"03", x"fa", x"03", x"fa", x"fe", x"fd",
    x"03", x"fa", x"02", x"ff", x"03", x"02", x"fd", x"03",
    x"03", x"04", x"01", x"03", x"03", x"f8", x"01", x"01",
    x"fe", x"ff", x"fc", x"fe", x"ff", x"02", x"ff", x"fc",
    x"03", x"fa", x"fd", x"ff", x"fa", x"fb", x"04", x"fc",
    x"ff", x"02", x"01", x"fb", x"00", x"fb", x"02", x"fe",
    x"fb", x"fb", x"ff", x"01", x"fc", x"fe", x"f8", x"fb",
    x"fe", x"03", x"fc", x"fc", x"ff", x"03", x"fb", x"f8",
    x"02", x"01", x"fe", x"f9", x"fe", x"fb", x"f9", x"01",
    x"01", x"fe", x"fe", x"fe", x"fd", x"00", x"00", x"02",
    x"fb", x"fe", x"ff", x"fe", x"fe", x"fd", x"fd", x"fd",
    x"03", x"fd", x"fb", x"02", x"00", x"01", x"fb", x"02",
    x"fb", x"fd", x"00", x"ff", x"fb", x"01", x"fe", x"00",
    x"01", x"ff", x"01", x"03", x"02", x"fa", x"02", x"fa",
    x"fe", x"01", x"fb", x"03", x"02", x"00", x"02", x"fb",
    x"fe", x"00", x"fd", x"fe", x"01", x"04", x"fb", x"fd",
    x"fd", x"fc", x"fd", x"fe", x"03", x"fe", x"00", x"03",
    x"fa", x"ff", x"04", x"fe", x"fb", x"fd", x"00", x"fe",
    x"ff", x"01", x"fa", x"fd", x"fb", x"fe", x"ff", x"01",
    x"fa", x"03", x"ff", x"ff", x"05", x"fe", x"fd", x"fb",
    x"fd", x"fb", x"02", x"f7", x"04", x"00", x"00", x"00",
    x"fa", x"fa", x"fd", x"fc", x"fd", x"f8", x"04", x"fe",
    x"00", x"ff", x"f7", x"f8", x"01", x"f8", x"fe", x"f6",
    x"fc", x"00", x"fa", x"fc", x"00", x"fa", x"01", x"fd",
    x"fc", x"fb", x"fd", x"fb", x"00", x"ff", x"fa", x"fc",
    x"fb", x"00", x"fc", x"fd", x"00", x"f7", x"f9", x"fe",
    x"00", x"fc", x"03", x"00", x"ff", x"fd", x"fa", x"f6",
    x"f7", x"fd", x"fd", x"f8", x"fa", x"fe", x"00", x"fd",
    x"03", x"01", x"01", x"fe", x"ff", x"04", x"01", x"fb",
    x"02", x"ff", x"fd", x"fe", x"fc", x"f7", x"fe", x"00",
    x"ff", x"fe", x"02", x"01", x"05", x"00", x"fc", x"fc",
    x"fb", x"fb", x"01", x"fb", x"f8", x"fa", x"fd", x"fc",
    x"fb", x"ff", x"fd", x"fa", x"fe", x"fb", x"fb", x"04",
    x"02", x"fe", x"fa", x"fe", x"ff", x"fc", x"ff", x"f9",
    x"02", x"fa", x"fd", x"fd", x"00", x"fb", x"fb", x"fe",
    x"fc", x"01", x"fd", x"01", x"01", x"04", x"f9", x"fb",
    x"fb", x"02", x"fc", x"fe", x"03", x"ff", x"00", x"fc",
    x"05", x"ff", x"00", x"ff", x"02", x"fd", x"fa", x"ff",
    x"00", x"fb", x"00", x"ff", x"f7", x"ff", x"00", x"fd",
    x"fc", x"03", x"02", x"fd", x"f8", x"00", x"fd", x"fb",
    x"03", x"01", x"fa", x"ff", x"fc", x"00", x"f9", x"f8",
    x"ff", x"ff", x"fd", x"fb", x"03", x"04", x"fc", x"fc",
    x"ff", x"00", x"f7", x"03", x"fe", x"04", x"fe", x"fa",
    x"01", x"fe", x"fb", x"fc", x"ff", x"fd", x"fc", x"fd",
    x"ff", x"fc", x"f8", x"03", x"03", x"f9", x"ff", x"fb",
    x"fe", x"f7", x"fe", x"f9", x"01", x"fd", x"f7", x"ff",
    x"fc", x"ff", x"ff", x"fd", x"f7", x"fa", x"00", x"04",
    x"fc", x"04", x"ff", x"04", x"fc", x"02", x"fb", x"fc",
    x"03", x"04", x"03", x"05", x"fe", x"fd", x"ff", x"fe",
    x"00", x"f7", x"fb", x"fe", x"fa", x"f6", x"01", x"ff",
    x"ff", x"00", x"ff", x"ff", x"fd", x"fa", x"f7", x"fc",
    x"fd", x"00", x"ff", x"03", x"fe", x"fe", x"fc", x"fc",
    x"f9", x"f9", x"f7", x"fd", x"00", x"04", x"02", x"fc",
    x"f8", x"03", x"01", x"04", x"fb", x"04", x"f7", x"fd",
    x"ff", x"fc", x"ff", x"fe", x"00", x"00", x"fc", x"fb",
    x"00", x"fd", x"00", x"fd", x"fe", x"fc", x"fe", x"fb",
    x"fb", x"fb", x"03", x"00", x"02", x"fa", x"ff", x"fe",
    x"fb", x"01", x"ff", x"03", x"05", x"fb", x"fa", x"ff",
    x"00", x"01", x"04", x"03", x"03", x"fe", x"01", x"01",
    x"f8", x"00", x"fd", x"ff", x"fd", x"f9", x"04", x"fe",
    x"f7", x"fa", x"fd", x"ff", x"04", x"fd", x"fd", x"01",
    x"02", x"02", x"fb", x"02", x"04", x"fd", x"01", x"03",
    x"fd", x"fc", x"fb", x"00", x"03", x"03", x"ff", x"fa",
    x"fc", x"02", x"f8", x"fd", x"f7", x"f9", x"fd", x"fd",
    x"fc", x"f9", x"04", x"fc", x"ff", x"02", x"f8", x"f8",
    x"ff", x"00", x"ff", x"ff", x"fd", x"fd", x"02", x"ff",
    x"fd", x"00", x"fd", x"fa", x"fb", x"00", x"01", x"f7",
    x"fe", x"03", x"00", x"fe", x"f9", x"04", x"00", x"fe",
    x"f8", x"f7", x"fd", x"f7", x"ff", x"fb", x"01", x"00",
    x"fc", x"00", x"fa", x"01", x"fe", x"00", x"f8", x"ff",
    x"f8", x"00", x"fa", x"fa", x"f8", x"fb", x"ff", x"02",
    x"fc", x"fb", x"04", x"00", x"02", x"00", x"03", x"fc",
    x"04", x"fe", x"00", x"04", x"fc", x"03", x"00", x"02",
    x"fe", x"fd", x"fe", x"00", x"f9", x"00", x"f9", x"04",
    x"f9", x"ff", x"05", x"00", x"f9", x"fe", x"f7", x"01",
    x"00", x"fc", x"03", x"04", x"fd", x"00", x"04", x"ff",
    x"fc", x"f9", x"fd", x"fb", x"02", x"ff", x"fa", x"ff",
    x"fd", x"ff", x"fd", x"ff", x"fb", x"ff", x"04", x"fb",
    x"04", x"fb", x"fe", x"05", x"fc", x"f8", x"f8", x"02",
    x"04", x"fb", x"01", x"fb", x"01", x"fd", x"fc", x"00",
    x"05", x"05", x"f8", x"01", x"04", x"f7", x"fd", x"fd",
    x"f7", x"fd", x"fa", x"fb", x"00", x"01", x"04", x"fd",
    x"00", x"fc", x"03", x"fa", x"f9", x"f8", x"fd", x"fe",
    x"fe", x"fe", x"fb", x"f9", x"00", x"ff", x"f7", x"f7",
    x"fd", x"00", x"02", x"fd", x"fc", x"fb", x"fc", x"00",
    x"fd", x"00", x"fa", x"01", x"05", x"fe", x"fd", x"f7",
    x"fe", x"f9", x"f9", x"fd", x"fe", x"ff", x"fe", x"fe",
    x"ff", x"ff", x"00", x"fb", x"01", x"f7", x"f9", x"fb",
    x"fd", x"f9", x"f8", x"03", x"ff", x"fc", x"04", x"ff",
    x"27", x"2c", x"f2", x"1f", x"22", x"e0", x"22", x"0d",
    x"e7", x"12", x"de", x"d3", x"9f", x"eb", x"ca", x"18",
    x"e1", x"dc", x"dc", x"01", x"f3", x"0e", x"e9", x"08",
    x"06", x"d2", x"1f", x"0c", x"02", x"45", x"16", x"11",
    x"1d", x"12", x"19", x"0f", x"e9", x"08", x"b5", x"1f",
    x"e9", x"f5", x"f7", x"ef", x"0a", x"b5", x"bc", x"c0",
    x"92", x"e3", x"b6", x"72", x"d7", x"bd", x"7f", x"34",
    x"21", x"14", x"f4", x"f7", x"23", x"ed", x"fd", x"bc",
    x"ef", x"f5", x"05", x"f9", x"18", x"06", x"23", x"13",
    x"f8", x"f9", x"07", x"e7", x"04", x"ff", x"eb", x"e8",
    x"ee", x"f0", x"cf", x"c3", x"9d", x"f1", x"f7", x"c0",
    x"e8", x"e5", x"62", x"29", x"1d", x"1b", x"0c", x"2a",
    x"f1", x"3b", x"3a", x"0f", x"e0", x"fb", x"e9", x"01",
    x"0e", x"1a", x"1c", x"1e", x"ce", x"de", x"a0", x"fd",
    x"73", x"6f", x"1a", x"94", x"7f", x"cd", x"da", x"8f",
    x"eb", x"e0", x"35", x"c9", x"c0", x"51", x"13", x"5a",
    x"9e", x"af", x"80", x"76", x"ea", x"c4", x"8c", x"02",
    x"26", x"0c", x"0e", x"1b", x"23", x"0b", x"09", x"0c",
    x"99", x"06", x"f2", x"09", x"dc", x"0b", x"e8", x"2e",
    x"19", x"ff", x"01", x"04", x"fe", x"fb", x"fe", x"fc",
    x"00", x"ff", x"ea", x"7d", x"c7", x"ad", x"69", x"af",
    x"02", x"ed", x"eb", x"d3", x"00", x"e6", x"9c", x"fa",
    x"c3", x"88", x"ae", x"7b", x"1b", x"1f", x"f2", x"f2",
    x"25", x"26", x"ef", x"24", x"1e", x"c9", x"b7", x"05",
    x"df", x"da", x"fa", x"fe", x"d6", x"b6", x"eb", x"fb",
    x"1a", x"02", x"0c", x"02", x"15", x"0f", x"ff", x"c6",
    x"f5", x"e1", x"e7", x"de", x"00", x"e3", x"fc", x"0d",
    x"df", x"25", x"24", x"b9", x"19", x"fd", x"c6", x"05",
    x"04", x"21", x"19", x"04", x"f7", x"28", x"1a", x"a1",
    x"3a", x"1f", x"eb", x"0e", x"02", x"e8", x"09", x"fa",
    x"b9", x"ab", x"78", x"04", x"fe", x"fa", x"01", x"fe",
    x"f9", x"fd", x"fa", x"01", x"dc", x"df", x"c2", x"fa",
    x"bb", x"c2", x"b8", x"d9", x"c2", x"2e", x"23", x"62",
    x"54", x"51", x"40", x"48", x"3d", x"2f", x"e7", x"e3",
    x"e4", x"d5", x"b5", x"df", x"1b", x"1d", x"12", x"ec",
    x"b0", x"cf", x"bf", x"72", x"92", x"a7", x"4d", x"5b",
    x"26", x"27", x"22", x"17", x"07", x"13", x"19", x"00",
    x"15", x"bc", x"0b", x"18", x"91", x"11", x"93", x"ff",
    x"24", x"c5", x"69", x"4d", x"39", x"24", x"0f", x"0f",
    x"0a", x"f6", x"0d", x"60", x"46", x"10", x"24", x"e5",
    x"bc", x"0a", x"da", x"e8", x"01", x"04", x"02", x"08",
    x"0d", x"13", x"0d", x"04", x"02", x"20", x"17", x"f9",
    x"16", x"09", x"f8", x"36", x"24", x"12", x"d9", x"16",
    x"13", x"28", x"fc", x"12", x"7a", x"0b", x"fd", x"b1",
    x"08", x"0b", x"26", x"13", x"09", x"04", x"04", x"04",
    x"fd", x"ff", x"fc", x"04", x"fe", x"fe", x"fc", x"fb",
    x"03", x"f6", x"f6", x"fa", x"b6", x"ba", x"e6", x"1f",
    x"c0", x"a2", x"ba", x"f9", x"0e", x"12", x"fa", x"14",
    x"e3", x"b2", x"7b", x"1e", x"f6", x"0a", x"bd", x"e0",
    x"dd", x"c2", x"ea", x"f6", x"f2", x"0e", x"22", x"bd",
    x"d0", x"e5", x"e6", x"e5", x"06", x"08", x"28", x"11",
    x"ef", x"ee", x"de", x"9d", x"c6", x"df", x"86", x"c1",
    x"e9", x"99", x"f0", x"1a", x"f3", x"04", x"f9", x"d0",
    x"af", x"e8", x"d5", x"9c", x"c5", x"e9", x"e2", x"b6",
    x"fe", x"00", x"fc", x"fe", x"05", x"fc", x"03", x"00",
    x"05", x"03", x"04", x"01", x"ff", x"fe", x"fc", x"00",
    x"fd", x"ff", x"d9", x"db", x"cf", x"22", x"f5", x"de",
    x"1c", x"2f", x"1c", x"1c", x"31", x"f5", x"fc", x"ff",
    x"a4", x"e8", x"0e", x"d1", x"d3", x"d0", x"99", x"c9",
    x"d8", x"b2", x"e5", x"0e", x"f4", x"db", x"cd", x"bf",
    x"fb", x"c7", x"e1", x"ea", x"a2", x"be", x"cd", x"f3",
    x"f9", x"2a", x"e0", x"03", x"c4", x"0d", x"13", x"9c",
    x"1f", x"0d", x"6b", x"18", x"0c", x"6d", x"02", x"04",
    x"04", x"1a", x"0e", x"17", x"1b", x"0b", x"f2", x"04",
    x"17", x"e6", x"e2", x"fb", x"f6", x"f5", x"0b", x"f3",
    x"13", x"fa", x"10", x"ee", x"df", x"19", x"1e", x"0b",
    x"13", x"0d", x"18", x"a8", x"71", x"6a", x"ba", x"cd",
    x"88", x"ef", x"dc", x"f9", x"0b", x"5e", x"44", x"1a",
    x"ed", x"d1", x"ee", x"03", x"11", x"f6", x"29", x"e4",
    x"fc", x"09", x"de", x"d9", x"f9", x"a6", x"da", x"3a",
    x"0f", x"ec", x"1e", x"2c", x"b9", x"1e", x"13", x"ca",
    x"14", x"2c", x"f3", x"06", x"23", x"e8", x"2f", x"34",
    x"3b", x"f9", x"b7", x"2f", x"10", x"f8", x"2e", x"38",
    x"32", x"0a", x"f3", x"0b", x"bf", x"db", x"ed", x"11",
    x"c7", x"da", x"1c", x"2f", x"26", x"17", x"01", x"18",
    x"f5", x"08", x"08", x"ff", x"d9", x"e5", x"f9", x"e3",
    x"05", x"e9", x"14", x"06", x"1f", x"b9", x"a7", x"ce",
    x"c2", x"bc", x"f6", x"e3", x"d3", x"94", x"f7", x"dd",
    x"c4", x"b0", x"b6", x"f6", x"ed", x"05", x"e8", x"30",
    x"27", x"f6", x"f2", x"07", x"27", x"f9", x"e2", x"cf",
    x"ab", x"6c", x"f9", x"e2", x"00", x"0c", x"ff", x"f3",
    x"a5", x"a1", x"8e", x"ec", x"af", x"de", x"0e", x"da",
    x"17", x"b5", x"a2", x"77", x"6b", x"80", x"c1", x"d1",
    x"aa", x"22", x"82", x"0d", x"20", x"4b", x"ec", x"f1",
    x"f9", x"d6", x"fb", x"36", x"31", x"1c", x"22", x"33",
    x"1d", x"3e", x"0b", x"1b", x"ff", x"ce", x"05", x"3f",
    x"f8", x"0e", x"3b", x"28", x"1a", x"a7", x"9c", x"32",
    x"05", x"c8", x"1d", x"29", x"09", x"26", x"fb", x"2f",
    x"24", x"e1", x"cd", x"ff", x"03", x"0e", x"19", x"c4",
    x"e3", x"e9", x"ae", x"eb", x"1f", x"e0", x"f2", x"30",
    x"da", x"1b", x"00", x"0e", x"0e", x"04", x"3f", x"f9",
    x"ba", x"04", x"fd", x"fc", x"04", x"ff", x"04", x"03",
    x"ff", x"05", x"b4", x"d6", x"c4", x"88", x"f2", x"0f",
    x"0d", x"27", x"0c", x"93", x"ac", x"96", x"8f", x"bc",
    x"cf", x"79", x"96", x"e1", x"2e", x"2c", x"fc", x"d6",
    x"07", x"d8", x"ca", x"08", x"ec", x"15", x"f0", x"ea",
    x"f8", x"fe", x"04", x"ff", x"08", x"07", x"40", x"24",
    x"13", x"10", x"17", x"22", x"f7", x"17", x"13", x"ee",
    x"d8", x"e5", x"d9", x"fd", x"fb", x"da", x"ec", x"d6",
    x"21", x"1e", x"0f", x"43", x"e4", x"fc", x"10", x"ca",
    x"ef", x"0f", x"24", x"30", x"33", x"09", x"0f", x"42",
    x"1e", x"eb", x"d8", x"c6", x"da", x"0b", x"00", x"f9",
    x"2d", x"1b", x"03", x"fe", x"02", x"fc", x"f9", x"05",
    x"01", x"01", x"fd", x"fc", x"9a", x"9f", x"cd", x"a1",
    x"da", x"f8", x"da", x"ee", x"f2", x"27", x"f9", x"38",
    x"38", x"29", x"01", x"44", x"2f", x"77", x"df", x"bf",
    x"16", x"cb", x"dc", x"14", x"08", x"d9", x"eb", x"9f",
    x"94", x"d1", x"d8", x"d3", x"d5", x"1e", x"08", x"12",
    x"d8", x"cf", x"fd", x"1b", x"3c", x"62", x"33", x"38",
    x"23", x"b8", x"b5", x"ea", x"73", x"80", x"05", x"d3",
    x"e5", x"05", x"14", x"5d", x"58", x"41", x"1e", x"48",
    x"23", x"34", x"33", x"dc", x"ef", x"ed", x"19", x"02",
    x"12", x"22", x"15", x"11", x"01", x"ff", x"05", x"f9",
    x"03", x"02", x"01", x"05", x"fe", x"d0", x"e5", x"e5",
    x"ef", x"f8", x"10", x"22", x"05", x"07", x"4c", x"e2",
    x"fb", x"29", x"03", x"04", x"4f", x"07", x"05", x"1d",
    x"09", x"03", x"2f", x"09", x"fc", x"34", x"1a", x"fb",
    x"03", x"01", x"01", x"fc", x"05", x"05", x"fe", x"fc",
    x"00", x"1b", x"c6", x"d4", x"6a", x"b9", x"b8", x"1c",
    x"f2", x"1c", x"4e", x"17", x"ca", x"38", x"fa", x"e8",
    x"32", x"10", x"f8", x"ed", x"0f", x"22", x"01", x"f7",
    x"f0", x"c8", x"f2", x"ec", x"7c", x"8d", x"d7", x"8e",
    x"ca", x"26", x"07", x"ef", x"1d", x"4c", x"2e", x"08",
    x"de", x"f3", x"e9", x"03", x"ee", x"ec", x"8a", x"f3",
    x"fb", x"b1", x"de", x"e7", x"ec", x"09", x"04", x"db",
    x"dd", x"14", x"d8", x"d7", x"e8", x"1a", x"00", x"0e",
    x"03", x"ff", x"f9", x"05", x"04", x"02", x"fd", x"00",
    x"05", x"f7", x"ff", x"ff", x"05", x"fb", x"ff", x"00",
    x"06", x"03", x"5f", x"38", x"0a", x"2e", x"31", x"05",
    x"33", x"1f", x"ee", x"35", x"2d", x"11", x"26", x"1c",
    x"0e", x"05", x"09", x"f1", x"a3", x"9b", x"c4", x"e1",
    x"9b", x"e4", x"2c", x"b3", x"a9", x"d8", x"f0", x"2c",
    x"25", x"24", x"33", x"14", x"45", x"40", x"18", x"08",
    x"12", x"c7", x"b8", x"00", x"fa", x"0b", x"1b", x"35",
    x"0c", x"11", x"4c", x"f9", x"fd", x"75", x"fa", x"f7",
    x"88", x"43", x"31", x"2a", x"1f", x"1e", x"22", x"bb",
    x"e5", x"06", x"f3", x"fa", x"10", x"db", x"d4", x"1a",
    x"ec", x"df", x"0a", x"02", x"06", x"11", x"15", x"2d",
    x"02", x"2d", x"1b", x"00", x"e7", x"bd", x"0d", x"12",
    x"f7", x"36", x"0b", x"1b", x"1d", x"04", x"ea", x"20",
    x"43", x"19", x"2a", x"1d", x"21", x"e7", x"ee", x"09",
    x"fd", x"f3", x"e5", x"fa", x"ee", x"dc", x"e4", x"3b",
    x"27", x"ee", x"0a", x"0b", x"4b", x"23", x"f6", x"47",
    x"53", x"50", x"2a", x"2a", x"3e", x"18", x"20", x"f1",
    x"eb", x"e4", x"cb", x"12", x"e2", x"1a", x"11", x"ea",
    x"e4", x"49", x"d7", x"de", x"25", x"0b", x"24", x"24",
    x"29", x"08", x"f1", x"e6", x"d9", x"d2", x"9c", x"95",
    x"be", x"d0", x"d6", x"10", x"f4", x"d4", x"fe", x"c7",
    x"f0", x"eb", x"10", x"1c", x"b2", x"94", x"df", x"b4",
    x"bb", x"f0", x"81", x"92", x"99", x"c8", x"16", x"42",
    x"93", x"1c", x"24", x"f8", x"28", x"10", x"6d", x"c6",
    x"ed", x"4d", x"08", x"f0", x"14", x"d6", x"01", x"54",
    x"ea", x"58", x"d9", x"46", x"41", x"3a", x"3c", x"0e",
    x"6a", x"df", x"f7", x"07", x"07", x"ff", x"08", x"f1",
    x"f5", x"e3", x"35", x"4a", x"d5", x"fc", x"f7", x"03",
    x"16", x"13", x"c9", x"11", x"0f", x"f9", x"ea", x"ee",
    x"33", x"da", x"0d", x"d0", x"09", x"f8", x"ed", x"02",
    x"fb", x"1d", x"13", x"e2", x"17", x"4f", x"36", x"4b",
    x"13", x"d1", x"3e", x"cf", x"c0", x"a8", x"9a", x"a0",
    x"cf", x"b7", x"f2", x"20", x"29", x"38", x"1c", x"22",
    x"09", x"c7", x"09", x"05", x"50", x"36", x"16", x"ae",
    x"c5", x"07", x"b2", x"c9", x"1e", x"b8", x"13", x"27",
    x"e6", x"28", x"4f", x"40", x"41", x"28", x"ec", x"d7",
    x"eb", x"01", x"01", x"ff", x"ff", x"00", x"fe", x"fa",
    x"fb", x"ff", x"b8", x"76", x"e9", x"a0", x"d7", x"65",
    x"16", x"23", x"36", x"ec", x"dc", x"d2", x"dc", x"de",
    x"fa", x"ce", x"0e", x"16", x"07", x"ee", x"c2", x"db",
    x"e4", x"12", x"19", x"21", x"11", x"c6", x"0b", x"01",
    x"00", x"e0", x"ed", x"ee", x"bc", x"ea", x"ca", x"1a",
    x"1f", x"2f", x"17", x"1c", x"fd", x"d3", x"c6", x"9f",
    x"de", x"fa", x"ba", x"e0", x"f4", x"d3", x"c8", x"b3",
    x"d5", x"98", x"e2", x"ed", x"b3", x"e3", x"18", x"1e",
    x"0e", x"0a", x"e3", x"ff", x"f8", x"f6", x"28", x"1e",
    x"1c", x"0a", x"ee", x"fc", x"05", x"fd", x"06", x"fc",
    x"fa", x"06", x"05", x"00", x"f9", x"fd", x"fb", x"f7",
    x"fc", x"f2", x"fc", x"fd", x"dd", x"1d", x"fc", x"f7",
    x"14", x"0d", x"f1", x"f7", x"26", x"01", x"fa", x"fd",
    x"3f", x"2d", x"e6", x"fd", x"a9", x"13", x"11", x"db",
    x"a9", x"df", x"2d", x"2e", x"31", x"1c", x"1b", x"7c",
    x"d5", x"d3", x"f3", x"f8", x"16", x"34", x"0f", x"0a",
    x"ee", x"2e", x"ed", x"f0", x"38", x"1c", x"1b", x"f6",
    x"28", x"d8", x"e4", x"38", x"e7", x"f4", x"27", x"02",
    x"fc", x"eb", x"8e", x"0e", x"01", x"e3", x"1e", x"01",
    x"39", x"4a", x"f1", x"e7", x"ad", x"ff", x"e3", x"b6",
    x"ee", x"33", x"25", x"1c", x"04", x"f9", x"f8", x"08",
    x"04", x"ff", x"02", x"05", x"05", x"ca", x"06", x"33",
    x"2a", x"03", x"1a", x"0b", x"0a", x"fe", x"fc", x"06",
    x"c4", x"fc", x"a7", x"d6", x"e9", x"fa", x"06", x"03",
    x"1f", x"01", x"e2", x"f7", x"ee", x"17", x"18", x"ee",
    x"fb", x"ff", x"fe", x"fa", x"00", x"02", x"fc", x"05",
    x"04", x"18", x"cd", x"79", x"c7", x"87", x"da", x"3c",
    x"18", x"22", x"f4", x"ac", x"80", x"d0", x"e6", x"f9",
    x"20", x"f1", x"0b", x"a4", x"e1", x"ae", x"ee", x"e9",
    x"17", x"19", x"27", x"00", x"d2", x"9e", x"a7", x"b2",
    x"ad", x"04", x"e3", x"f1", x"0a", x"e5", x"38", x"11",
    x"c1", x"f1", x"0b", x"23", x"0e", x"fb", x"ff", x"40",
    x"0b", x"77", x"93", x"ef", x"b4", x"d5", x"1a", x"c2",
    x"fe", x"28", x"c9", x"db", x"f4", x"d4", x"05", x"0f",
    x"07", x"f9", x"fb", x"03", x"f9", x"ff", x"fa", x"06",
    x"ff", x"fe", x"f9", x"fb", x"01", x"f9", x"fa", x"fd",
    x"fa", x"ff", x"12", x"0f", x"3e", x"02", x"f8", x"e8",
    x"a6", x"a9", x"8d", x"31", x"5f", x"13", x"24", x"06",
    x"31", x"1f", x"08", x"17", x"d8", x"de", x"22", x"d5",
    x"f6", x"fd", x"b4", x"d6", x"0c", x"dc", x"36", x"20",
    x"1c", x"fc", x"14", x"d2", x"fb", x"34", x"db", x"df",
    x"f1", x"2b", x"bd", x"ec", x"a8", x"e4", x"22", x"f5",
    x"dc", x"f7", x"47", x"c5", x"d9", x"4c", x"0d", x"10",
    x"1d", x"16", x"d3", x"eb", x"07", x"c4", x"c7", x"c8",
    x"e1", x"d6", x"19", x"1d", x"61", x"08", x"30", x"0d",
    x"df", x"dd", x"b1", x"0b", x"fc", x"ee", x"f5", x"19",
    x"fe", x"2a", x"21", x"12", x"1a", x"22", x"01", x"03",
    x"f2", x"40", x"21", x"d2", x"ee", x"2a", x"1c", x"09",
    x"2f", x"03", x"14", x"fd", x"f4", x"f0", x"44", x"2e",
    x"12", x"39", x"17", x"e5", x"ff", x"12", x"e3", x"04",
    x"f3", x"34", x"1c", x"fc", x"4d", x"26", x"f4", x"d1",
    x"17", x"00", x"d2", x"e7", x"1e", x"35", x"2e", x"03",
    x"0f", x"1d", x"1f", x"fd", x"f0", x"23", x"14", x"3b",
    x"3b", x"32", x"01", x"04", x"c1", x"dd", x"ea", x"0e",
    x"0e", x"05", x"32", x"53", x"44", x"1a", x"37", x"2c",
    x"ed", x"14", x"1a", x"db", x"20", x"24", x"09", x"e2",
    x"f0", x"f4", x"d2", x"ee", x"17", x"24", x"1c", x"e3",
    x"09", x"29", x"fa", x"06", x"20", x"36", x"14", x"9d",
    x"47", x"17", x"c7", x"f8", x"27", x"25", x"ec", x"d7",
    x"ec", x"27", x"f2", x"fd", x"21", x"e3", x"f7", x"b9",
    x"a9", x"09", x"84", x"68", x"d6", x"ca", x"de", x"26",
    x"b0", x"aa", x"c6", x"b6", x"b1", x"cb", x"dd", x"06",
    x"2d", x"f9", x"1b", x"da", x"d1", x"02", x"36", x"ff",
    x"38", x"42", x"44", x"3f", x"20", x"28", x"43", x"26",
    x"1b", x"fd", x"2c", x"e6", x"14", x"fb", x"d9", x"0c",
    x"0f", x"0b", x"1c", x"0e", x"d1", x"ed", x"02", x"fa",
    x"03", x"f9", x"12", x"ee", x"f2", x"0d", x"13", x"f6",
    x"06", x"12", x"31", x"fd", x"0a", x"36", x"48", x"27",
    x"2d", x"f8", x"e8", x"f8", x"d2", x"ee", x"fa", x"6e",
    x"3b", x"0c", x"17", x"05", x"18", x"eb", x"f2", x"07",
    x"e5", x"da", x"bf", x"ef", x"00", x"9f", x"c5", x"c7",
    x"f4", x"01", x"fe", x"fd", x"fc", x"04", x"03", x"00",
    x"fd", x"02", x"89", x"32", x"2c", x"fa", x"a1", x"c6",
    x"07", x"f6", x"ef", x"03", x"05", x"b0", x"1c", x"0f",
    x"d9", x"35", x"18", x"17", x"4a", x"36", x"b8", x"f3",
    x"0e", x"f4", x"34", x"d4", x"f0", x"32", x"20", x"15",
    x"2f", x"28", x"31", x"cf", x"b9", x"d5", x"3b", x"0d",
    x"01", x"2a", x"15", x"16", x"da", x"e5", x"f6", x"cd",
    x"bd", x"a1", x"c6", x"e5", x"ce", x"e9", x"cc", x"05",
    x"e6", x"dc", x"0b", x"12", x"c1", x"12", x"31", x"0c",
    x"14", x"19", x"20", x"28", x"14", x"04", x"fe", x"2b",
    x"f5", x"02", x"08", x"f5", x"19", x"11", x"07", x"1a",
    x"e9", x"eb", x"c2", x"f7", x"f4", x"fa", x"fa", x"03",
    x"fa", x"fb", x"fb", x"fa", x"fa", x"9d", x"c1", x"b4",
    x"da", x"cd", x"98", x"ce", x"b5", x"18", x"44", x"1d",
    x"18", x"1c", x"ef", x"38", x"25", x"14", x"2e", x"03",
    x"15", x"14", x"11", x"2a", x"fb", x"fb", x"12", x"9d",
    x"b3", x"9a", x"bf", x"bd", x"91", x"fe", x"e5", x"17",
    x"e2", x"2a", x"03", x"ea", x"04", x"10", x"1d", x"d4",
    x"f8", x"0a", x"f9", x"07", x"de", x"e8", x"07", x"0a",
    x"17", x"33", x"0a", x"41", x"1d", x"fc", x"d4", x"f8",
    x"14", x"ee", x"b6", x"d4", x"f7", x"ad", x"cd", x"e1",
    x"c2", x"ff", x"24", x"00", x"01", x"0e", x"0a", x"03",
    x"03", x"10", x"08", x"fb", x"10", x"6b", x"16", x"23",
    x"ec", x"0b", x"0b", x"23", x"0e", x"06", x"53", x"ff",
    x"42", x"45", x"ff", x"19", x"49", x"2e", x"22", x"c4",
    x"b9", x"f1", x"34", x"fa", x"0e", x"49", x"2a", x"24",
    x"04", x"fd", x"fb", x"fe", x"01", x"04", x"fb", x"03",
    x"fd", x"11", x"df", x"e9", x"0c", x"e8", x"fc", x"c7",
    x"03", x"0d", x"c9", x"65", x"94", x"aa", x"7f", x"bc",
    x"cd", x"cf", x"d5", x"14", x"0a", x"31", x"f1", x"ed",
    x"12", x"f3", x"04", x"1d", x"0f", x"3d", x"37", x"0a",
    x"05", x"1c", x"fd", x"03", x"ff", x"e3", x"f3", x"d8",
    x"d7", x"d5", x"d5", x"d7", x"09", x"1b", x"71", x"00",
    x"eb", x"05", x"ec", x"be", x"08", x"08", x"d0", x"2f",
    x"36", x"29", x"1e", x"1f", x"15", x"16", x"04", x"fd",
    x"fe", x"00", x"00", x"fb", x"fe", x"06", x"fc", x"fe",
    x"00", x"02", x"01", x"01", x"fc", x"ff", x"fd", x"fe",
    x"02", x"00", x"32", x"3e", x"02", x"29", x"1f", x"fd",
    x"2e", x"1a", x"fa", x"1e", x"fc", x"41", x"2f", x"f9",
    x"25", x"2d", x"df", x"f2", x"3a", x"62", x"5b", x"35",
    x"43", x"2a", x"10", x"24", x"1c", x"d0", x"ea", x"ef",
    x"d1", x"c4", x"e1", x"13", x"44", x"fc", x"de", x"fa",
    x"07", x"dc", x"e0", x"d0", x"eb", x"fc", x"ea", x"04",
    x"d9", x"ce", x"2b", x"ef", x"fa", x"28", x"09", x"fc",
    x"5c", x"fc", x"3f", x"40", x"2d", x"14", x"35", x"26",
    x"fa", x"ae", x"db", x"1f", x"60", x"16", x"e4", x"2b",
    x"12", x"f3", x"61", x"f1", x"1a", x"41", x"53", x"42",
    x"01", x"58", x"37", x"2f", x"f1", x"23", x"06", x"03",
    x"07", x"06", x"d4", x"cd", x"14", x"a9", x"ca", x"d8",
    x"c9", x"bf", x"39", x"3e", x"24", x"ed", x"f0", x"e8",
    x"f8", x"d8", x"cf", x"ad", x"e8", x"ec", x"e8", x"d2",
    x"27", x"80", x"c6", x"0e", x"04", x"da", x"1b", x"f7",
    x"b6", x"fe", x"15", x"ab", x"d3", x"1c", x"fb", x"db",
    x"e3", x"0f", x"6c", x"c0", x"f2", x"24", x"e7", x"1d",
    x"3d", x"b0", x"e9", x"03", x"15", x"df", x"0c", x"00",
    x"f7", x"d9", x"e0", x"d7", x"04", x"09", x"f0", x"e2",
    x"57", x"22", x"03", x"ff", x"0d", x"e9", x"f4", x"04",
    x"24", x"ee", x"d7", x"eb", x"26", x"f6", x"1c", x"bd",
    x"b8", x"e8", x"a0", x"a7", x"cf", x"ca", x"aa", x"fd",
    x"a9", x"b6", x"bd", x"1b", x"dc", x"15", x"cf", x"f1",
    x"d7", x"c6", x"ca", x"16", x"05", x"3d", x"47", x"f7",
    x"10", x"29", x"09", x"1d", x"d5", x"e4", x"cb", x"a8",
    x"0e", x"0c", x"28", x"e0", x"0f", x"ec", x"ad", x"a2",
    x"e7", x"c7", x"b9", x"10", x"1e", x"38", x"37", x"ff",
    x"61", x"6f", x"22", x"2a", x"fd", x"be", x"01", x"13",
    x"2f", x"e0", x"48", x"bb", x"f1", x"19", x"1a", x"35",
    x"3b", x"2d", x"72", x"60", x"1d", x"e9", x"e5", x"9e",
    x"d3", x"e2", x"a1", x"e3", x"cd", x"4d", x"12", x"18",
    x"f9", x"18", x"33", x"ef", x"01", x"3c", x"e3", x"dd",
    x"0e", x"28", x"20", x"04", x"03", x"04", x"15", x"7e",
    x"e8", x"b7", x"ed", x"0b", x"2f", x"3b", x"2b", x"38",
    x"a1", x"cf", x"58", x"b3", x"fb", x"51", x"f0", x"f0",
    x"e5", x"fb", x"fd", x"fb", x"05", x"fe", x"fb", x"00",
    x"05", x"00", x"13", x"1c", x"3f", x"54", x"1a", x"15",
    x"d9", x"f1", x"fc", x"f0", x"02", x"2c", x"0f", x"f2",
    x"23", x"32", x"45", x"bb", x"dc", x"fb", x"e4", x"dd",
    x"e3", x"ef", x"f6", x"f4", x"e8", x"01", x"fe", x"f1",
    x"f0", x"fc", x"e6", x"ef", x"b8", x"a0", x"1e", x"13",
    x"0c", x"f8", x"03", x"2b", x"ec", x"d7", x"f3", x"3d",
    x"1e", x"eb", x"f2", x"fa", x"f6", x"9a", x"ca", x"f0",
    x"41", x"51", x"3a", x"b4", x"0e", x"15", x"36", x"fc",
    x"17", x"18", x"f1", x"f7", x"f5", x"dd", x"ec", x"16",
    x"d6", x"7a", x"28", x"14", x"1a", x"d9", x"e6", x"f8",
    x"d2", x"c6", x"d3", x"0a", x"07", x"00", x"07", x"05",
    x"05", x"0c", x"0a", x"02", x"25", x"eb", x"ff", x"01",
    x"0f", x"fd", x"08", x"f1", x"24", x"08", x"17", x"19",
    x"e2", x"d4", x"cc", x"fb", x"19", x"3e", x"33", x"1e",
    x"04", x"ff", x"3d", x"34", x"13", x"13", x"ea", x"07",
    x"ff", x"00", x"14", x"12", x"01", x"e2", x"11", x"1a",
    x"0b", x"10", x"ef", x"c5", x"f4", x"ff", x"b6", x"d0",
    x"d4", x"e1", x"e4", x"16", x"ef", x"24", x"ee", x"d3",
    x"2e", x"1d", x"88", x"db", x"da", x"9d", x"c9", x"f6",
    x"aa", x"d8", x"f2", x"0b", x"23", x"11", x"fa", x"37",
    x"03", x"ae", x"3c", x"24", x"0f", x"00", x"02", x"09",
    x"0c", x"10", x"ff", x"fd", x"fd", x"21", x"e6", x"f2",
    x"d9", x"cf", x"02", x"f0", x"0f", x"12", x"f5", x"1c",
    x"08", x"e1", x"1e", x"09", x"aa", x"0f", x"fe", x"e1",
    x"e1", x"0e", x"c0", x"e0", x"f0", x"19", x"fd", x"fe",
    x"02", x"fe", x"ff", x"03", x"ff", x"03", x"00", x"00",
    x"03", x"31", x"2d", x"38", x"08", x"23", x"31", x"10",
    x"20", x"22", x"47", x"1c", x"0a", x"3c", x"38", x"34",
    x"14", x"d5", x"f1", x"26", x"23", x"15", x"fd", x"2e",
    x"29", x"e3", x"15", x"2f", x"13", x"27", x"e1", x"d6",
    x"d7", x"da", x"e5", x"ca", x"af", x"19", x"21", x"10",
    x"2b", x"2b", x"28", x"ba", x"d4", x"d7", x"f4", x"c2",
    x"f4", x"fa", x"d5", x"d7", x"ee", x"f5", x"02", x"25",
    x"ff", x"e8", x"23", x"f8", x"cc", x"ee", x"07", x"0f",
    x"fa", x"01", x"01", x"00", x"05", x"03", x"03", x"08",
    x"01", x"03", x"01", x"00", x"ff", x"08", x"05", x"ff",
    x"08", x"fe", x"ad", x"d4", x"fe", x"ae", x"9c", x"b6",
    x"d6", x"b1", x"e2", x"08", x"ef", x"00", x"fb", x"01",
    x"0a", x"ff", x"e7", x"e1", x"fa", x"e1", x"f4", x"a0",
    x"9e", x"b6", x"e9", x"d3", x"45", x"e8", x"02", x"e0",
    x"07", x"06", x"d4", x"d7", x"e8", x"ac", x"f8", x"21",
    x"db", x"25", x"f1", x"e1", x"1d", x"2f", x"08", x"ef",
    x"ed", x"08", x"a8", x"c3", x"f7", x"19", x"15", x"18",
    x"c5", x"b1", x"0c", x"ef", x"02", x"31", x"73", x"dc",
    x"03", x"3b", x"f4", x"f0", x"23", x"28", x"2e", x"28",
    x"14", x"2d", x"d4", x"b0", x"b3", x"ca", x"a3", x"af",
    x"2f", x"05", x"f2", x"e3", x"e3", x"eb", x"16", x"c9",
    x"c7", x"a8", x"ac", x"bd", x"1f", x"4a", x"f9", x"2c",
    x"21", x"05", x"26", x"20", x"2a", x"ed", x"0a", x"55",
    x"e0", x"df", x"fc", x"01", x"ef", x"fc", x"de", x"55",
    x"32", x"94", x"05", x"20", x"cb", x"f6", x"cd", x"ce",
    x"ff", x"d8", x"c1", x"d9", x"c5", x"67", x"d1", x"32",
    x"fd", x"fe", x"f8", x"03", x"f5", x"fb", x"fb", x"fa",
    x"fb", x"04", x"01", x"fa", x"02", x"ff", x"fe", x"fc",
    x"fd", x"f9", x"fd", x"f8", x"fb", x"fa", x"01", x"00",
    x"02", x"00", x"fe", x"fc", x"f7", x"f8", x"fd", x"01",
    x"f9", x"f9", x"f9", x"fa", x"fe", x"fd", x"fd", x"04",
    x"f8", x"fb", x"02", x"04", x"f9", x"fa", x"fd", x"03",
    x"fd", x"fe", x"fc", x"fd", x"fa", x"ff", x"fe", x"f8",
    x"fe", x"04", x"03", x"f5", x"fd", x"01", x"fb", x"03",
    x"fd", x"fd", x"04", x"00", x"01", x"03", x"f7", x"fb",
    x"fd", x"f9", x"ff", x"fb", x"fb", x"fa", x"02", x"fd",
    x"fd", x"03", x"fe", x"f9", x"fc", x"fa", x"fc", x"f8",
    x"fa", x"01", x"fe", x"03", x"fc", x"04", x"fd", x"fc",
    x"fe", x"01", x"f9", x"04", x"03", x"ff", x"fc", x"f9",
    x"f5", x"fc", x"fa", x"fe", x"00", x"05", x"06", x"03",
    x"fa", x"01", x"02", x"05", x"ff", x"fc", x"01", x"01",
    x"fb", x"fd", x"ff", x"01", x"fb", x"fc", x"02", x"fd",
    x"fb", x"00", x"05", x"ff", x"fc", x"fd", x"fc", x"fa",
    x"fb", x"04", x"01", x"fe", x"03", x"f9", x"fe", x"f8",
    x"fe", x"fe", x"02", x"01", x"03", x"f5", x"fb", x"03",
    x"fe", x"02", x"01", x"03", x"03", x"04", x"00", x"ff",
    x"fd", x"fd", x"fe", x"fb", x"04", x"ff", x"fd", x"01",
    x"fd", x"fa", x"fe", x"fc", x"02", x"00", x"00", x"ff",
    x"fe", x"fd", x"f8", x"ff", x"02", x"fc", x"02", x"03",
    x"fa", x"01", x"ff", x"fc", x"f8", x"fc", x"03", x"fb",
    x"fa", x"00", x"ff", x"f8", x"f8", x"fc", x"01", x"fc",
    x"fb", x"fb", x"f8", x"fd", x"ff", x"01", x"ff", x"01",
    x"01", x"fb", x"ff", x"fd", x"fd", x"00", x"fb", x"ff",
    x"fe", x"fd", x"fd", x"fc", x"f9", x"fa", x"f5", x"fe",
    x"fd", x"fb", x"04", x"ff", x"05", x"f8", x"fe", x"ff",
    x"fd", x"f6", x"fb", x"fa", x"03", x"02", x"fa", x"fd",
    x"f9", x"f9", x"02", x"fe", x"04", x"02", x"02", x"ff",
    x"04", x"02", x"01", x"fe", x"fc", x"ff", x"f9", x"fd",
    x"f9", x"f9", x"fd", x"fe", x"f9", x"fc", x"01", x"01",
    x"04", x"f9", x"ff", x"fd", x"01", x"02", x"fc", x"fa",
    x"00", x"03", x"00", x"fc", x"fc", x"fb", x"fa", x"fb",
    x"03", x"00", x"03", x"00", x"00", x"ff", x"f8", x"f5",
    x"fc", x"f9", x"01", x"fc", x"02", x"fe", x"fb", x"ff",
    x"00", x"04", x"06", x"fd", x"fd", x"07", x"f8", x"00",
    x"fe", x"ff", x"ff", x"ff", x"fc", x"f9", x"ff", x"00",
    x"f5", x"f5", x"fe", x"02", x"ff", x"04", x"fe", x"03",
    x"02", x"f6", x"fe", x"fa", x"04", x"00", x"ff", x"fc",
    x"fc", x"06", x"02", x"ff", x"02", x"ff", x"fb", x"fc",
    x"01", x"01", x"ff", x"01", x"fc", x"f9", x"05", x"00",
    x"fd", x"f9", x"fe", x"00", x"fc", x"05", x"ff", x"ff",
    x"fe", x"01", x"fd", x"ff", x"fc", x"fc", x"ff", x"fc",
    x"fe", x"00", x"05", x"05", x"03", x"05", x"04", x"ff",
    x"fe", x"fd", x"01", x"fd", x"fd", x"00", x"fe", x"fd",
    x"fc", x"f8", x"ff", x"fa", x"01", x"03", x"fd", x"02",
    x"02", x"04", x"fc", x"02", x"00", x"fb", x"06", x"fa",
    x"fe", x"01", x"fa", x"fd", x"03", x"fb", x"03", x"fd",
    x"01", x"fa", x"fd", x"fe", x"00", x"06", x"fb", x"01",
    x"fb", x"fe", x"ff", x"01", x"fb", x"fa", x"ff", x"fa",
    x"00", x"fe", x"06", x"01", x"03", x"fd", x"02", x"fd",
    x"fc", x"02", x"fd", x"fe", x"f9", x"fb", x"ff", x"ff",
    x"fb", x"ff", x"fb", x"02", x"00", x"04", x"ff", x"fb",
    x"01", x"05", x"00", x"ff", x"fd", x"fa", x"fe", x"02",
    x"fd", x"05", x"ff", x"fa", x"fd", x"ff", x"fc", x"fe",
    x"ff", x"f6", x"fe", x"01", x"fc", x"00", x"02", x"00",
    x"00", x"fe", x"ff", x"fd", x"04", x"02", x"01", x"fd",
    x"ff", x"ff", x"fe", x"fb", x"05", x"02", x"fc", x"fc",
    x"00", x"fb", x"fd", x"f8", x"f8", x"f7", x"05", x"fb",
    x"02", x"06", x"f9", x"ff", x"02", x"fd", x"fb", x"f9",
    x"fc", x"01", x"00", x"ff", x"f7", x"fd", x"ff", x"00",
    x"fe", x"02", x"fd", x"ff", x"fb", x"ff", x"fe", x"03",
    x"f9", x"ff", x"fe", x"fa", x"01", x"fb", x"fd", x"f8",
    x"f5", x"ff", x"04", x"f9", x"03", x"01", x"fc", x"01",
    x"fb", x"fa", x"f7", x"05", x"02", x"ff", x"fc", x"fd",
    x"01", x"00", x"f8", x"00", x"fb", x"00", x"00", x"04",
    x"01", x"fc", x"ff", x"fd", x"fc", x"fe", x"f9", x"01",
    x"fd", x"03", x"ff", x"fb", x"ff", x"00", x"fd", x"04",
    x"00", x"01", x"fc", x"fd", x"f9", x"01", x"01", x"fb",
    x"f9", x"ff", x"fd", x"fe", x"01", x"00", x"f9", x"fa",
    x"e4", x"12", x"62", x"d9", x"fb", x"4a", x"10", x"1e",
    x"1c", x"12", x"09", x"bf", x"f3", x"fa", x"1a", x"e4",
    x"2b", x"2e", x"28", x"30", x"6e", x"49", x"41", x"23",
    x"29", x"16", x"db", x"ca", x"c1", x"e7", x"f9", x"1d",
    x"14", x"e9", x"c0", x"0f", x"11", x"51", x"17", x"31",
    x"3a", x"d9", x"31", x"c9", x"ab", x"f6", x"c9", x"f6",
    x"e1", x"fb", x"1a", x"fc", x"38", x"f2", x"e0", x"e9",
    x"d3", x"00", x"25", x"00", x"1a", x"2b", x"da", x"0e",
    x"e9", x"e3", x"f6", x"eb", x"15", x"0b", x"0e", x"11",
    x"11", x"1f", x"30", x"08", x"f5", x"cb", x"07", x"ce",
    x"b6", x"fd", x"09", x"0b", x"01", x"f7", x"b5", x"06",
    x"ec", x"bb", x"8a", x"46", x"f2", x"01", x"42", x"d6",
    x"3d", x"20", x"fe", x"bc", x"ef", x"1b", x"9d", x"2c",
    x"19", x"9f", x"21", x"06", x"e6", x"2b", x"41", x"f9",
    x"1e", x"42", x"24", x"3f", x"23", x"2f", x"57", x"62",
    x"13", x"03", x"d4", x"01", x"13", x"25", x"d8", x"c1",
    x"c5", x"f1", x"e6", x"f5", x"e7", x"de", x"ca", x"fa",
    x"09", x"34", x"0b", x"1b", x"08", x"df", x"a6", x"d7",
    x"db", x"bb", x"9d", x"d8", x"bc", x"ec", x"17", x"f3",
    x"15", x"01", x"03", x"ff", x"fc", x"01", x"ff", x"01",
    x"02", x"01", x"bd", x"2c", x"00", x"b0", x"e5", x"e4",
    x"f7", x"04", x"14", x"24", x"49", x"23", x"02", x"d5",
    x"a6", x"fe", x"de", x"ac", x"ec", x"42", x"38", x"1c",
    x"1b", x"bd", x"06", x"fc", x"0b", x"1c", x"ee", x"fe",
    x"46", x"23", x"17", x"25", x"de", x"c7", x"ff", x"c4",
    x"f7", x"d8", x"d8", x"1d", x"3a", x"68", x"28", x"2c",
    x"26", x"3f", x"3d", x"2b", x"17", x"27", x"29", x"10",
    x"27", x"1d", x"2f", x"ae", x"23", x"21", x"6f", x"1d",
    x"14", x"05", x"22", x"e0", x"db", x"01", x"e2", x"dc",
    x"f6", x"16", x"30", x"19", x"e6", x"2f", x"10", x"fd",
    x"03", x"fc", x"17", x"fa", x"01", x"f9", x"0c", x"fe",
    x"fb", x"07", x"02", x"01", x"18", x"e9", x"f6", x"05",
    x"f9", x"f5", x"e4", x"d4", x"dc", x"0a", x"a8", x"bc",
    x"0b", x"d6", x"d3", x"2d", x"d1", x"e5", x"1d", x"1a",
    x"30", x"f2", x"f8", x"fb", x"0c", x"fb", x"e7", x"1f",
    x"1e", x"01", x"0f", x"ff", x"c4", x"11", x"c7", x"a9",
    x"da", x"ff", x"08", x"f2", x"0f", x"0b", x"e1", x"f8",
    x"0d", x"01", x"17", x"fd", x"05", x"23", x"d9", x"fe",
    x"f3", x"f7", x"a4", x"95", x"a8", x"a3", x"b0", x"dc",
    x"c2", x"05", x"df", x"5f", x"36", x"2b", x"27", x"05",
    x"eb", x"0b", x"e4", x"c2", x"01", x"f9", x"0e", x"fe",
    x"f8", x"fc", x"fe", x"fc", x"04", x"52", x"2c", x"19",
    x"21", x"fc", x"ab", x"0a", x"d3", x"e8", x"07", x"72",
    x"40", x"f6", x"1e", x"26", x"0b", x"1a", x"00", x"0c",
    x"22", x"16", x"d7", x"fd", x"f7", x"f6", x"18", x"fc",
    x"02", x"fe", x"fe", x"00", x"ff", x"fd", x"05", x"fd",
    x"fe", x"28", x"25", x"4d", x"03", x"03", x"19", x"04",
    x"d2", x"bb", x"07", x"2c", x"2b", x"0f", x"49", x"01",
    x"f3", x"f0", x"c4", x"49", x"1b", x"1d", x"1b", x"f4",
    x"dd", x"22", x"fa", x"f0", x"47", x"43", x"7a", x"04",
    x"28", x"e8", x"fd", x"09", x"3e", x"1e", x"52", x"5d",
    x"2c", x"39", x"24", x"2b", x"16", x"e6", x"4a", x"f1",
    x"e3", x"ce", x"fc", x"27", x"fc", x"da", x"1c", x"23",
    x"46", x"c6", x"13", x"d0", x"ef", x"fe", x"ef", x"f1",
    x"00", x"05", x"04", x"09", x"fb", x"02", x"02", x"03",
    x"02", x"06", x"05", x"fc", x"02", x"03", x"09", x"fe",
    x"ff", x"fd", x"e9", x"c9", x"da", x"c8", x"ea", x"13",
    x"08", x"1c", x"fc", x"cd", x"e6", x"30", x"f2", x"eb",
    x"e1", x"1f", x"0a", x"b5", x"2d", x"26", x"f7", x"21",
    x"fa", x"e9", x"05", x"fb", x"11", x"ea", x"eb", x"d8",
    x"fe", x"00", x"f3", x"f7", x"b4", x"dd", x"43", x"e4",
    x"ee", x"fc", x"0b", x"08", x"c5", x"0c", x"1b", x"0c",
    x"d5", x"01", x"d4", x"21", x"21", x"fc", x"29", x"0e",
    x"91", x"dd", x"34", x"8c", x"1d", x"3a", x"19", x"2d",
    x"38", x"33", x"e1", x"c9", x"e3", x"ef", x"03", x"f7",
    x"09", x"17", x"cb", x"9d", x"05", x"0f", x"f0", x"21",
    x"12", x"16", x"f9", x"d3", x"fc", x"c5", x"ba", x"e7",
    x"3a", x"03", x"16", x"ff", x"30", x"f4", x"f9", x"fe",
    x"ce", x"00", x"f9", x"f5", x"ef", x"30", x"0a", x"ef",
    x"1c", x"db", x"17", x"2f", x"fe", x"16", x"cb", x"86",
    x"b7", x"de", x"f4", x"21", x"de", x"0b", x"ff", x"f1",
    x"94", x"8d", x"fd", x"c0", x"da", x"1a", x"0e", x"d1",
    x"d6", x"d9", x"b7", x"fc", x"08", x"19", x"30", x"03",
    x"d9", x"e4", x"28", x"18", x"1b", x"06", x"25", x"11",
    x"eb", x"e7", x"c3", x"f0", x"0a", x"fc", x"13", x"fb",
    x"c5", x"dc", x"f6", x"09", x"d7", x"ef", x"f9", x"24",
    x"16", x"e9", x"ea", x"dd", x"c3", x"ef", x"f3", x"fd",
    x"17", x"2a", x"15", x"e8", x"c0", x"f2", x"ff", x"db",
    x"f6", x"01", x"e1", x"46", x"f9", x"f5", x"f8", x"14",
    x"1d", x"34", x"06", x"16", x"e8", x"cc", x"fa", x"c3",
    x"d8", x"e8", x"b7", x"ca", x"b5", x"37", x"47", x"57",
    x"b1", x"af", x"5a", x"b1", x"b3", x"c9", x"01", x"22",
    x"62", x"e5", x"01", x"ea", x"8a", x"ea", x"c5", x"ab",
    x"eb", x"16", x"28", x"fb", x"ff", x"0f", x"30", x"16",
    x"13", x"d7", x"f6", x"1e", x"03", x"0d", x"33", x"0b",
    x"05", x"72", x"07", x"d6", x"01", x"8e", x"b8", x"31",
    x"14", x"00", x"fe", x"ce", x"d1", x"a0", x"56", x"7e",
    x"ec", x"e8", x"e3", x"07", x"f8", x"47", x"e8", x"28",
    x"f0", x"b8", x"b2", x"c9", x"e5", x"e2", x"04", x"ee",
    x"17", x"20", x"dd", x"ea", x"fe", x"8e", x"c8", x"fc",
    x"33", x"0e", x"f4", x"3e", x"19", x"f7", x"cf", x"d0",
    x"07", x"02", x"00", x"fd", x"04", x"fd", x"02", x"ff",
    x"01", x"fd", x"d1", x"c0", x"0b", x"ad", x"81", x"b1",
    x"0b", x"30", x"1a", x"f3", x"f3", x"d8", x"f9", x"0d",
    x"f3", x"1e", x"ec", x"f6", x"b0", x"dc", x"b9", x"e3",
    x"d5", x"0e", x"25", x"01", x"f4", x"14", x"05", x"f2",
    x"20", x"12", x"00", x"6c", x"28", x"17", x"2a", x"0c",
    x"f6", x"f1", x"08", x"06", x"f3", x"c0", x"2e", x"98",
    x"09", x"e5", x"f2", x"1f", x"16", x"db", x"f7", x"17",
    x"0f", x"33", x"ec", x"2c", x"dc", x"06", x"32", x"b8",
    x"0d", x"dc", x"cd", x"e9", x"ef", x"1e", x"5a", x"16",
    x"dc", x"c8", x"cc", x"f2", x"e9", x"ee", x"01", x"24",
    x"2c", x"18", x"35", x"06", x"05", x"ff", x"05", x"fc",
    x"fc", x"fe", x"f5", x"fb", x"a8", x"d6", x"cc", x"d6",
    x"b0", x"c0", x"fd", x"22", x"39", x"3b", x"e5", x"9f",
    x"28", x"25", x"20", x"4d", x"0d", x"eb", x"be", x"c8",
    x"fe", x"e6", x"d7", x"eb", x"a7", x"b8", x"dc", x"cf",
    x"ba", x"96", x"c5", x"c6", x"db", x"0a", x"f6", x"1c",
    x"80", x"92", x"d8", x"fa", x"f5", x"f2", x"23", x"36",
    x"27", x"f4", x"0b", x"07", x"fe", x"f8", x"22", x"d9",
    x"d1", x"24", x"fd", x"00", x"de", x"21", x"00", x"08",
    x"2a", x"0d", x"04", x"ac", x"d1", x"b7", x"ff", x"f1",
    x"06", x"75", x"49", x"19", x"02", x"f7", x"04", x"fb",
    x"02", x"f7", x"01", x"fe", x"04", x"e1", x"c9", x"fa",
    x"9d", x"1d", x"23", x"b1", x"fd", x"fd", x"21", x"b8",
    x"8a", x"4a", x"9d", x"af", x"ca", x"bc", x"f0", x"31",
    x"56", x"10", x"16", x"e9", x"fd", x"d8", x"de", x"d3",
    x"fe", x"02", x"02", x"03", x"04", x"03", x"05", x"01",
    x"01", x"e5", x"e2", x"f1", x"fa", x"f2", x"ea", x"f1",
    x"00", x"07", x"ca", x"aa", x"a6", x"ca", x"c7", x"bf",
    x"32", x"25", x"1b", x"04", x"e0", x"d0", x"0d", x"25",
    x"26", x"20", x"07", x"e7", x"eb", x"08", x"33", x"95",
    x"ed", x"23", x"ce", x"cc", x"ec", x"bf", x"ba", x"0d",
    x"34", x"5b", x"34", x"12", x"0e", x"04", x"f6", x"11",
    x"1c", x"cf", x"e2", x"6e", x"bb", x"04", x"12", x"c2",
    x"dc", x"1b", x"dc", x"f1", x"01", x"f5", x"d7", x"ed",
    x"04", x"04", x"fe", x"01", x"fe", x"04", x"01", x"01",
    x"02", x"00", x"fd", x"05", x"fd", x"fd", x"fc", x"fd",
    x"00", x"fd", x"06", x"03", x"fd", x"0c", x"16", x"e6",
    x"01", x"fc", x"df", x"1a", x"08", x"b3", x"2a", x"f6",
    x"02", x"30", x"1f", x"43", x"c5", x"eb", x"d9", x"24",
    x"3b", x"fa", x"36", x"4e", x"2d", x"d7", x"fd", x"cc",
    x"03", x"f6", x"fe", x"61", x"23", x"2c", x"0c", x"0e",
    x"09", x"d2", x"ea", x"23", x"5b", x"50", x"9e", x"03",
    x"1d", x"f6", x"7b", x"2d", x"fb", x"54", x"ff", x"f3",
    x"11", x"1a", x"0c", x"23", x"1d", x"d7", x"69", x"d3",
    x"0c", x"16", x"c2", x"d9", x"41", x"49", x"20", x"4b",
    x"54", x"fb", x"e5", x"0e", x"fe", x"22", x"f3", x"d8",
    x"15", x"09", x"29", x"14", x"22", x"0e", x"bc", x"ef",
    x"f2", x"ff", x"10", x"1d", x"c8", x"be", x"9c", x"d5",
    x"a4", x"a0", x"51", x"08", x"2c", x"ed", x"f8", x"fa",
    x"41", x"1b", x"db", x"08", x"f9", x"0b", x"ff", x"f8",
    x"ad", x"0f", x"ee", x"e1", x"0c", x"e9", x"ed", x"18",
    x"1f", x"fc", x"37", x"43", x"2d", x"64", x"1a", x"f7",
    x"fe", x"1c", x"19", x"18", x"3c", x"40", x"28", x"35",
    x"ef", x"3b", x"f7", x"e8", x"62", x"0f", x"fc", x"19",
    x"1c", x"f7", x"0f", x"0f", x"e0", x"f8", x"e0", x"b4",
    x"12", x"d2", x"c9", x"ff", x"1c", x"24", x"e3", x"e4",
    x"39", x"f6", x"e5", x"04", x"de", x"09", x"9a", x"d2",
    x"e6", x"b0", x"f1", x"da", x"05", x"2a", x"35", x"cd",
    x"e7", x"4b", x"1b", x"f5", x"38", x"e2", x"f8", x"10",
    x"1c", x"e6", x"ee", x"2a", x"17", x"14", x"f9", x"ed",
    x"7b", x"21", x"07", x"21", x"fb", x"05", x"08", x"ef",
    x"0c", x"fa", x"e2", x"df", x"f8", x"f5", x"f9", x"00",
    x"66", x"f3", x"f9", x"ea", x"c7", x"b2", x"0b", x"22",
    x"fc", x"ae", x"50", x"31", x"bc", x"0b", x"22", x"c5",
    x"38", x"15", x"f5", x"ea", x"00", x"27", x"ed", x"01",
    x"27", x"23", x"28", x"12", x"1f", x"07", x"35", x"f5",
    x"0e", x"0a", x"f3", x"02", x"e2", x"f0", x"c9", x"d4",
    x"08", x"b9", x"da", x"e8", x"b3", x"cd", x"11", x"02",
    x"c8", x"9c", x"a7", x"b2", x"a2", x"c4", x"ec", x"ea",
    x"dc", x"e8", x"d5", x"d4", x"fb", x"12", x"e9", x"cc",
    x"f3", x"e8", x"fd", x"1f", x"33", x"f9", x"fe", x"10",
    x"5f", x"ff", x"04", x"fd", x"03", x"01", x"fd", x"03",
    x"03", x"fd", x"ee", x"c6", x"df", x"e9", x"be", x"c7",
    x"f7", x"f3", x"1e", x"11", x"d2", x"92", x"1b", x"12",
    x"cd", x"1e", x"35", x"2a", x"2c", x"fb", x"ef", x"16",
    x"d0", x"94", x"e7", x"18", x"00", x"03", x"a5", x"80",
    x"f4", x"d8", x"f4", x"f0", x"12", x"53", x"f0", x"0f",
    x"0b", x"16", x"1d", x"e4", x"2d", x"41", x"28", x"09",
    x"ce", x"b2", x"1e", x"da", x"fc", x"fe", x"18", x"28",
    x"10", x"fc", x"2e", x"07", x"21", x"ed", x"d4", x"29",
    x"ec", x"3a", x"ed", x"ba", x"25", x"06", x"d3", x"e7",
    x"1f", x"43", x"f4", x"f7", x"e5", x"ad", x"f4", x"49",
    x"c1", x"1e", x"57", x"fb", x"fc", x"05", x"fe", x"02",
    x"fb", x"03", x"fc", x"fd", x"cb", x"8a", x"de", x"ee",
    x"a6", x"af", x"f4", x"c6", x"ad", x"11", x"19", x"22",
    x"06", x"26", x"0d", x"03", x"01", x"0e", x"1b", x"12",
    x"0b", x"eb", x"a3", x"e3", x"13", x"0a", x"e3", x"fa",
    x"c6", x"06", x"e0", x"f7", x"e6", x"02", x"e8", x"ff",
    x"fd", x"f2", x"f2", x"eb", x"eb", x"c5", x"f5", x"df",
    x"75", x"e1", x"d2", x"c2", x"dc", x"01", x"fd", x"0a",
    x"ea", x"0e", x"e7", x"19", x"2b", x"17", x"fa", x"25",
    x"14", x"f5", x"02", x"e3", x"1c", x"0d", x"28", x"0f",
    x"09", x"05", x"f6", x"f2", x"0a", x"05", x"03", x"09",
    x"02", x"09", x"09", x"01", x"06", x"15", x"c1", x"7a",
    x"3f", x"a1", x"a1", x"ff", x"b2", x"a8", x"41", x"1f",
    x"fb", x"f5", x"b6", x"b2", x"ff", x"c1", x"cf", x"fd",
    x"27", x"19", x"e7", x"21", x"c9", x"ec", x"d4", x"c7",
    x"03", x"03", x"ff", x"00", x"fe", x"ff", x"03", x"01",
    x"fb", x"50", x"ff", x"0e", x"28", x"db", x"04", x"52",
    x"05", x"c3", x"0a", x"d3", x"f0", x"08", x"df", x"11",
    x"35", x"17", x"0a", x"04", x"14", x"29", x"49", x"f5",
    x"3c", x"19", x"1c", x"3a", x"1d", x"58", x"3e", x"3a",
    x"bd", x"0a", x"f9", x"d8", x"bf", x"04", x"3e", x"4c",
    x"f2", x"27", x"3c", x"08", x"37", x"1d", x"0a", x"19",
    x"06", x"fa", x"03", x"0d", x"34", x"01", x"fa", x"c7",
    x"03", x"df", x"df", x"ec", x"3e", x"f4", x"f4", x"13",
    x"05", x"01", x"fe", x"ff", x"fc", x"fb", x"fb", x"05",
    x"03", x"fd", x"fd", x"fd", x"04", x"00", x"01", x"fa",
    x"fb", x"01", x"2e", x"b7", x"c8", x"ec", x"19", x"19",
    x"0c", x"fa", x"32", x"d7", x"2e", x"0b", x"0e", x"29",
    x"9d", x"f3", x"d9", x"9c", x"e1", x"e6", x"bb", x"ee",
    x"0f", x"35", x"ed", x"dd", x"1c", x"e0", x"bd", x"e1",
    x"f2", x"d4", x"f0", x"29", x"fb", x"ec", x"f5", x"17",
    x"07", x"b0", x"07", x"e3", x"12", x"21", x"35", x"ea",
    x"f3", x"3b", x"18", x"1c", x"34", x"2d", x"07", x"14",
    x"34", x"fa", x"f8", x"4b", x"20", x"e6", x"50", x"f7",
    x"de", x"e4", x"fe", x"33", x"e2", x"15", x"45", x"fe",
    x"28", x"1f", x"15", x"f5", x"2a", x"21", x"f6", x"13",
    x"fb", x"fe", x"bb", x"11", x"ee", x"e0", x"22", x"fb",
    x"eb", x"1a", x"c2", x"e8", x"ef", x"1c", x"35", x"08",
    x"fe", x"1e", x"3e", x"1a", x"33", x"1e", x"12", x"10",
    x"19", x"21", x"01", x"11", x"db", x"bd", x"19", x"43",
    x"3c", x"1d", x"fd", x"f5", x"12", x"10", x"b6", x"f3",
    x"0f", x"46", x"16", x"06", x"3c", x"c8", x"f1", x"1c",
    x"fb", x"00", x"fd", x"00", x"fb", x"ff", x"fb", x"fe",
    x"02", x"03", x"fc", x"00", x"02", x"fd", x"04", x"fc",
    x"ff", x"03", x"fe", x"03", x"03", x"fc", x"fe", x"fe",
    x"04", x"fd", x"fb", x"00", x"fd", x"fb", x"f6", x"fa",
    x"fc", x"fd", x"ff", x"ff", x"fd", x"fb", x"02", x"fe",
    x"fc", x"fc", x"03", x"fe", x"f8", x"ff", x"fc", x"fd",
    x"ff", x"fc", x"01", x"00", x"fd", x"fe", x"fb", x"fc",
    x"03", x"fb", x"fc", x"fd", x"01", x"00", x"ff", x"00",
    x"04", x"fd", x"fd", x"fe", x"01", x"fd", x"04", x"00",
    x"fa", x"fb", x"fe", x"03", x"fc", x"ff", x"fb", x"fb",
    x"00", x"fe", x"ff", x"ff", x"fe", x"fc", x"fa", x"03",
    x"fd", x"01", x"fe", x"fc", x"fd", x"fa", x"03", x"02",
    x"00", x"fe", x"01", x"fb", x"fa", x"f3", x"01", x"fd",
    x"f8", x"fc", x"02", x"02", x"03", x"fd", x"ff", x"fb",
    x"fc", x"fb", x"ff", x"ff", x"ff", x"fc", x"00", x"02",
    x"fc", x"fe", x"03", x"fc", x"fe", x"f9", x"fd", x"fd",
    x"03", x"fb", x"fb", x"05", x"03", x"01", x"f6", x"fc",
    x"03", x"00", x"fc", x"fc", x"fb", x"01", x"fb", x"fb",
    x"02", x"fa", x"03", x"02", x"fb", x"f8", x"fa", x"ff",
    x"fc", x"05", x"fc", x"03", x"fe", x"fd", x"fd", x"ff",
    x"fc", x"fe", x"ff", x"fa", x"fc", x"fe", x"fc", x"01",
    x"fa", x"fe", x"fe", x"03", x"fc", x"03", x"03", x"fa",
    x"02", x"fd", x"f9", x"fd", x"fe", x"00", x"ff", x"ff",
    x"05", x"04", x"fe", x"f8", x"02", x"03", x"01", x"fd",
    x"fd", x"fe", x"ff", x"fa", x"f8", x"00", x"fe", x"03",
    x"01", x"fa", x"02", x"ff", x"02", x"ff", x"00", x"01",
    x"fe", x"ff", x"00", x"04", x"ff", x"fc", x"ff", x"f9",
    x"04", x"03", x"fb", x"03", x"02", x"f8", x"04", x"fe",
    x"ff", x"fe", x"00", x"01", x"01", x"fa", x"01", x"04",
    x"fb", x"fb", x"ff", x"02", x"fd", x"fb", x"ff", x"ff",
    x"02", x"fd", x"03", x"fd", x"04", x"fc", x"fb", x"fe",
    x"02", x"ff", x"fd", x"fc", x"ff", x"fe", x"fd", x"00",
    x"fc", x"01", x"02", x"fe", x"f9", x"00", x"fd", x"ff",
    x"00", x"fa", x"fd", x"ff", x"fc", x"fe", x"fc", x"03",
    x"fa", x"fd", x"fe", x"f7", x"fd", x"fa", x"fd", x"03",
    x"01", x"00", x"fb", x"fd", x"02", x"fb", x"fb", x"fa",
    x"02", x"fb", x"fb", x"f9", x"f9", x"00", x"f9", x"fd",
    x"fe", x"02", x"fb", x"f8", x"fa", x"fc", x"02", x"fc",
    x"00", x"02", x"ff", x"fd", x"00", x"03", x"fa", x"fc",
    x"fb", x"00", x"fc", x"ff", x"fd", x"ff", x"01", x"fb",
    x"f6", x"fc", x"fa", x"03", x"fb", x"00", x"fb", x"fc",
    x"03", x"fb", x"ff", x"04", x"01", x"fb", x"fc", x"fd",
    x"fe", x"03", x"02", x"fe", x"fe", x"fd", x"03", x"04",
    x"fd", x"01", x"fc", x"00", x"05", x"02", x"02", x"f9",
    x"03", x"00", x"fb", x"fc", x"02", x"03", x"fd", x"fd",
    x"04", x"fc", x"04", x"fc", x"02", x"fb", x"fc", x"fd",
    x"fd", x"03", x"00", x"01", x"03", x"00", x"fb", x"fd",
    x"01", x"01", x"fc", x"03", x"fb", x"fa", x"fb", x"fb",
    x"fc", x"fe", x"01", x"01", x"ff", x"02", x"fd", x"fd",
    x"fb", x"fe", x"02", x"ff", x"ff", x"00", x"fe", x"02",
    x"01", x"fb", x"fb", x"fd", x"02", x"ff", x"04", x"fb",
    x"fb", x"fe", x"fe", x"02", x"fe", x"f7", x"03", x"03",
    x"fd", x"02", x"03", x"01", x"fb", x"00", x"00", x"02",
    x"ff", x"fb", x"ff", x"fd", x"01", x"00", x"fa", x"ff",
    x"ff", x"fb", x"fc", x"03", x"04", x"fc", x"fc", x"fd",
    x"02", x"ff", x"02", x"fc", x"fd", x"00", x"fa", x"fe",
    x"ff", x"ff", x"01", x"fd", x"00", x"fc", x"fa", x"ff",
    x"01", x"f9", x"f8", x"fa", x"fa", x"00", x"fc", x"fc",
    x"fd", x"01", x"04", x"02", x"01", x"fa", x"fb", x"01",
    x"03", x"fc", x"01", x"00", x"00", x"03", x"fc", x"f9",
    x"fa", x"00", x"fd", x"fc", x"ff", x"fd", x"03", x"01",
    x"ff", x"fc", x"02", x"01", x"ff", x"03", x"fe", x"02",
    x"fd", x"fc", x"fd", x"00", x"01", x"ff", x"02", x"01",
    x"03", x"ff", x"02", x"fb", x"fe", x"01", x"00", x"03",
    x"fa", x"02", x"01", x"00", x"00", x"01", x"fe", x"03",
    x"04", x"fe", x"03", x"fd", x"00", x"fb", x"01", x"f8",
    x"fc", x"fa", x"fb", x"fe", x"03", x"fb", x"fa", x"fa",
    x"fc", x"ff", x"00", x"ff", x"00", x"fd", x"04", x"fa",
    x"fa", x"fb", x"fe", x"03", x"01", x"ff", x"fb", x"f9",
    x"fa", x"02", x"fc", x"00", x"02", x"fd", x"ff", x"00",
    x"ff", x"fd", x"fc", x"04", x"02", x"fe", x"00", x"02",
    x"01", x"fb", x"04", x"04", x"fd", x"fa", x"02", x"02",
    x"09", x"d8", x"bd", x"df", x"e4", x"f5", x"e3", x"f4",
    x"2d", x"db", x"0b", x"2a", x"e4", x"ce", x"ac", x"af",
    x"bc", x"e8", x"d8", x"07", x"1f", x"dd", x"f5", x"fd",
    x"04", x"03", x"12", x"d5", x"a0", x"cd", x"d5", x"f4",
    x"07", x"0f", x"11", x"c9", x"f2", x"ee", x"03", x"eb",
    x"d0", x"ce", x"f1", x"11", x"f5", x"fe", x"1d", x"0f",
    x"13", x"e4", x"11", x"cb", x"e9", x"dc", x"1e", x"15",
    x"dd", x"1c", x"37", x"13", x"1c", x"2e", x"20", x"1c",
    x"f7", x"28", x"23", x"1c", x"04", x"ef", x"c3", x"dd",
    x"ce", x"15", x"4e", x"18", x"31", x"29", x"f6", x"07",
    x"f1", x"1a", x"fc", x"e7", x"fb", x"c7", x"b9", x"cb",
    x"d3", x"b9", x"2d", x"21", x"14", x"ee", x"2d", x"07",
    x"f7", x"30", x"09", x"45", x"18", x"fa", x"47", x"13",
    x"0c", x"cf", x"30", x"18", x"35", x"cd", x"ec", x"c7",
    x"d0", x"ec", x"05", x"36", x"25", x"0c", x"21", x"38",
    x"09", x"31", x"26", x"fb", x"f4", x"86", x"02", x"f8",
    x"f9", x"32", x"24", x"22", x"38", x"1a", x"1d", x"1c",
    x"0a", x"08", x"de", x"db", x"f1", x"13", x"e7", x"f8",
    x"ec", x"10", x"26", x"06", x"23", x"1d", x"12", x"fe",
    x"1f", x"06", x"03", x"01", x"00", x"ff", x"fd", x"01",
    x"03", x"05", x"29", x"47", x"25", x"15", x"09", x"f7",
    x"df", x"fb", x"15", x"11", x"0e", x"fc", x"ff", x"cd",
    x"fa", x"6a", x"6d", x"f9", x"49", x"29", x"ee", x"37",
    x"e1", x"c7", x"b2", x"e3", x"0a", x"fa", x"ec", x"e9",
    x"da", x"e5", x"01", x"e0", x"c2", x"cc", x"ee", x"c5",
    x"cc", x"ea", x"d8", x"03", x"f7", x"23", x"1d", x"20",
    x"04", x"fd", x"0f", x"c9", x"e0", x"7d", x"7b", x"b5",
    x"35", x"28", x"25", x"0e", x"ec", x"07", x"df", x"2a",
    x"18", x"0c", x"05", x"0a", x"19", x"c1", x"f0", x"77",
    x"f7", x"ff", x"fd", x"21", x"30", x"fc", x"2c", x"ca",
    x"de", x"cb", x"bd", x"ff", x"fb", x"06", x"fe", x"f8",
    x"06", x"03", x"ff", x"0b", x"22", x"2a", x"03", x"15",
    x"07", x"df", x"23", x"aa", x"7a", x"12", x"19", x"09",
    x"01", x"c6", x"b6", x"2d", x"12", x"34", x"f6", x"f3",
    x"ef", x"1e", x"00", x"f5", x"40", x"4a", x"41", x"02",
    x"fd", x"20", x"18", x"0e", x"34", x"b0", x"87", x"92",
    x"fe", x"e1", x"1b", x"1d", x"2b", x"44", x"e5", x"06",
    x"10", x"25", x"31", x"14", x"f7", x"08", x"4b", x"dd",
    x"e1", x"82", x"66", x"0a", x"33", x"68", x"25", x"20",
    x"9f", x"fb", x"f3", x"19", x"f8", x"fa", x"d8", x"c7",
    x"f1", x"22", x"72", x"5d", x"fc", x"0d", x"08", x"fa",
    x"fd", x"f9", x"f9", x"fb", x"fd", x"22", x"f1", x"fe",
    x"d1", x"11", x"1e", x"f6", x"ec", x"d2", x"ea", x"e5",
    x"d6", x"b7", x"11", x"1c", x"f9", x"20", x"1f", x"0e",
    x"b0", x"d5", x"f0", x"24", x"4b", x"1e", x"27", x"37",
    x"f9", x"fc", x"01", x"03", x"ff", x"02", x"01", x"fd",
    x"00", x"f4", x"0a", x"fb", x"f6", x"f4", x"ef", x"36",
    x"fe", x"26", x"1e", x"47", x"22", x"23", x"2d", x"36",
    x"ef", x"ae", x"a7", x"f8", x"0c", x"1a", x"30", x"fb",
    x"d8", x"02", x"80", x"74", x"bd", x"f8", x"ed", x"ff",
    x"0f", x"34", x"15", x"02", x"f0", x"f0", x"fa", x"f7",
    x"f5", x"d9", x"fa", x"00", x"ed", x"ec", x"0d", x"fa",
    x"78", x"e3", x"e5", x"e9", x"f1", x"04", x"04", x"2a",
    x"44", x"23", x"16", x"ee", x"10", x"f2", x"f5", x"24",
    x"06", x"fe", x"09", x"02", x"08", x"fc", x"08", x"fd",
    x"01", x"ff", x"06", x"03", x"fb", x"ff", x"02", x"fc",
    x"03", x"01", x"01", x"0f", x"1a", x"f6", x"07", x"0d",
    x"05", x"f0", x"f5", x"17", x"46", x"45", x"0e", x"13",
    x"33", x"0d", x"12", x"04", x"05", x"05", x"ec", x"0a",
    x"10", x"d7", x"d0", x"e3", x"ef", x"20", x"38", x"24",
    x"37", x"42", x"0f", x"dc", x"ce", x"dc", x"f0", x"eb",
    x"ff", x"2d", x"48", x"0d", x"17", x"fe", x"ea", x"3e",
    x"2b", x"2c", x"21", x"17", x"0f", x"4c", x"46", x"41",
    x"f9", x"e8", x"ea", x"8f", x"99", x"df", x"c5", x"16",
    x"ea", x"dd", x"08", x"1d", x"f1", x"b2", x"86", x"f7",
    x"b7", x"bb", x"f5", x"e2", x"f0", x"e6", x"e8", x"1a",
    x"fd", x"f8", x"ef", x"1c", x"0f", x"f9", x"33", x"0d",
    x"05", x"8b", x"9a", x"12", x"07", x"30", x"03", x"d5",
    x"d5", x"f1", x"b0", x"96", x"b2", x"f4", x"0f", x"f2",
    x"0c", x"7d", x"92", x"ea", x"b7", x"71", x"1c", x"f7",
    x"ed", x"1c", x"00", x"fe", x"d7", x"15", x"23", x"e1",
    x"1d", x"40", x"d9", x"04", x"ff", x"cd", x"ef", x"b4"
  );

  type fc1_bias_128_t is array (0 to 127) of std_logic_vector(7 downto 0);
  constant fc1_bias : fc1_bias_128_t := (
    x"ff", x"ee", x"db", x"ff", x"f7", x"fc", x"0b", x"e3",
    x"f3", x"de", x"bb", x"e2", x"10", x"cd", x"d7", x"e6",
    x"c6", x"ea", x"f6", x"0c", x"f9", x"0f", x"e5", x"dc",
    x"f8", x"e4", x"e7", x"e9", x"ed", x"cd", x"d4", x"f5",
    x"11", x"e0", x"f9", x"f2", x"fe", x"fc", x"d8", x"f5",
    x"c6", x"ef", x"c6", x"ca", x"0a", x"f8", x"fe", x"e3",
    x"1d", x"f7", x"0a", x"e4", x"f9", x"21", x"02", x"fb",
    x"f2", x"eb", x"ee", x"df", x"07", x"f8", x"c9", x"f7",
    x"fd", x"e4", x"d9", x"e8", x"fb", x"e8", x"f9", x"de",
    x"f9", x"e3", x"f8", x"d7", x"07", x"d4", x"e7", x"ec",
    x"f0", x"00", x"f6", x"e9", x"fa", x"b6", x"f7", x"f6",
    x"04", x"f9", x"e1", x"e9", x"fe", x"03", x"ff", x"eb",
    x"06", x"fd", x"0a", x"e5", x"0b", x"fd", x"fc", x"f7",
    x"db", x"f0", x"eb", x"d8", x"03", x"ec", x"ec", x"f5",
    x"da", x"02", x"ff", x"fd", x"f9", x"0b", x"0a", x"f4",
    x"e8", x"f4", x"f7", x"dc", x"fb", x"f8", x"fa", x"c9"
  );

  type fc1_activation_post_process_eps_1_t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant fc1_activation_post_process_eps : fc1_activation_post_process_eps_1_t := (
    x"00"
  );

  type fc1_activation_post_process_min_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant fc1_activation_post_process_min_val : fc1_activation_post_process_min_val__t := (
    x"7b"
  );

  type fc1_activation_post_process_max_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant fc1_activation_post_process_max_val : fc1_activation_post_process_max_val__t := (
    x"99"
  );

  type fc2_weight_10_128_t is array (0 to 1279) of std_logic_vector(7 downto 0);
  constant fc2_weight : fc2_weight_10_128_t := (
    x"0f", x"df", x"0e", x"f7", x"fa", x"f8", x"cf", x"d6",
    x"f4", x"e2", x"df", x"14", x"1a", x"db", x"d2", x"dc",
    x"0c", x"14", x"d7", x"17", x"fb", x"06", x"d9", x"0c",
    x"04", x"07", x"ca", x"eb", x"14", x"ce", x"0b", x"06",
    x"c6", x"ba", x"ea", x"a8", x"06", x"16", x"0f", x"1a",
    x"c7", x"12", x"16", x"07", x"15", x"f7", x"03", x"09",
    x"de", x"f7", x"24", x"11", x"c9", x"12", x"b2", x"f2",
    x"ef", x"c1", x"bd", x"0b", x"e4", x"b8", x"0d", x"b2",
    x"fa", x"0c", x"08", x"da", x"e0", x"0d", x"f6", x"10",
    x"e5", x"0f", x"f9", x"0b", x"f7", x"c7", x"02", x"ba",
    x"01", x"fb", x"05", x"db", x"c3", x"16", x"16", x"11",
    x"c2", x"ee", x"a9", x"0b", x"02", x"be", x"ff", x"1d",
    x"18", x"00", x"b8", x"ff", x"23", x"c6", x"00", x"04",
    x"be", x"b7", x"e1", x"f5", x"da", x"0a", x"18", x"ff",
    x"da", x"b3", x"01", x"01", x"ff", x"c1", x"16", x"18",
    x"1a", x"cf", x"f3", x"e3", x"0f", x"cf", x"f7", x"d5",
    x"0a", x"09", x"fe", x"06", x"fe", x"0c", x"ae", x"c9",
    x"fb", x"cc", x"f5", x"14", x"f8", x"20", x"02", x"cc",
    x"f5", x"ff", x"03", x"fd", x"f6", x"93", x"f4", x"9b",
    x"f4", x"b1", x"ff", x"ef", x"a2", x"1b", x"14", x"ff",
    x"ec", x"0c", x"91", x"16", x"f4", x"0e", x"cc", x"a8",
    x"fa", x"05", x"05", x"01", x"1c", x"05", x"fd", x"d8",
    x"05", x"f1", x"1b", x"f4", x"8b", x"de", x"15", x"03",
    x"05", x"16", x"f4", x"8c", x"03", x"07", x"ba", x"d4",
    x"f8", x"b7", x"02", x"d3", x"ec", x"b3", x"ff", x"9e",
    x"00", x"0c", x"ff", x"fc", x"ba", x"16", x"0d", x"0b",
    x"fc", x"0a", x"0c", x"af", x"0c", x"e0", x"18", x"16",
    x"0b", x"0a", x"13", x"d3", x"fe", x"10", x"03", x"09",
    x"04", x"fb", x"b8", x"98", x"0f", x"a4", x"f5", x"05",
    x"04", x"c4", x"08", x"dc", x"15", x"99", x"05", x"c1",
    x"fa", x"10", x"fe", x"03", x"00", x"0f", x"08", x"7a",
    x"0a", x"02", x"01", x"06", x"c2", x"f3", x"f8", x"c0",
    x"d4", x"18", x"12", x"04", x"02", x"00", x"e3", x"02",
    x"04", x"0f", x"0c", x"07", x"e0", x"12", x"1a", x"16",
    x"27", x"0d", x"c8", x"d0", x"01", x"ec", x"0f", x"07",
    x"f8", x"08", x"d3", x"0c", x"17", x"13", x"08", x"07",
    x"b6", x"d0", x"f0", x"e0", x"ff", x"cf", x"f0", x"d3",
    x"f7", x"e1", x"13", x"09", x"d9", x"ff", x"f9", x"16",
    x"ec", x"f6", x"be", x"dc", x"c3", x"b3", x"13", x"fe",
    x"c6", x"16", x"d0", x"09", x"e8", x"e3", x"f3", x"01",
    x"04", x"08", x"0c", x"14", x"f3", x"cd", x"fc", x"ed",
    x"c6", x"c7", x"04", x"11", x"e3", x"10", x"e7", x"1f",
    x"c5", x"c2", x"0c", x"fe", x"0c", x"16", x"0e", x"dc",
    x"e6", x"ff", x"db", x"0f", x"fd", x"d8", x"f2", x"f3",
    x"c6", x"06", x"ef", x"02", x"d8", x"e5", x"f7", x"04",
    x"cc", x"d0", x"0e", x"0a", x"e8", x"09", x"cf", x"cc",
    x"08", x"c1", x"fc", x"09", x"f9", x"c7", x"eb", x"d3",
    x"07", x"e2", x"05", x"0d", x"f4", x"06", x"f5", x"ea",
    x"e2", x"e0", x"16", x"03", x"fb", x"09", x"e5", x"0a",
    x"02", x"15", x"e3", x"fe", x"d7", x"0e", x"0e", x"de",
    x"cf", x"0a", x"0b", x"0f", x"fd", x"16", x"f5", x"cf",
    x"f8", x"f8", x"0b", x"0c", x"d0", x"0e", x"09", x"02",
    x"dc", x"14", x"12", x"d8", x"02", x"cf", x"10", x"1d",
    x"1c", x"e3", x"d3", x"01", x"ea", x"ff", x"fa", x"14",
    x"f5", x"03", x"c7", x"0d", x"ed", x"cf", x"b4", x"f9",
    x"d4", x"10", x"11", x"0a", x"14", x"0a", x"df", x"d4",
    x"00", x"d9", x"06", x"b5", x"a6", x"10", x"fa", x"dc",
    x"10", x"f0", x"fc", x"c9", x"fe", x"e2", x"d7", x"f3",
    x"da", x"ee", x"db", x"e2", x"e2", x"f6", x"e2", x"ec",
    x"1a", x"ed", x"f2", x"0b", x"03", x"db", x"05", x"bd",
    x"e5", x"01", x"eb", x"ed", x"e2", x"12", x"fb", x"03",
    x"05", x"de", x"0a", x"1c", x"0f", x"04", x"f0", x"c1",
    x"0f", x"ca", x"03", x"fe", x"0a", x"fb", x"ed", x"eb",
    x"0f", x"0f", x"05", x"06", x"d5", x"e5", x"f8", x"d2",
    x"d2", x"10", x"d5", x"05", x"f7", x"06", x"0f", x"d2",
    x"f9", x"cc", x"07", x"0c", x"b1", x"c1", x"e8", x"f2",
    x"13", x"e2", x"0b", x"d6", x"f4", x"ca", x"14", x"13",
    x"04", x"cd", x"10", x"e8", x"15", x"0f", x"03", x"05",
    x"00", x"bc", x"11", x"db", x"fd", x"0e", x"e5", x"c3",
    x"06", x"06", x"db", x"06", x"e0", x"09", x"04", x"ed",
    x"c9", x"03", x"09", x"09", x"08", x"aa", x"ba", x"f2",
    x"d8", x"10", x"10", x"ca", x"e7", x"12", x"e2", x"0d",
    x"07", x"11", x"c3", x"0c", x"f3", x"df", x"f9", x"0e",
    x"e4", x"11", x"04", x"0d", x"ed", x"13", x"0c", x"b9",
    x"f0", x"09", x"08", x"de", x"fb", x"f2", x"cf", x"0a",
    x"ac", x"0b", x"16", x"b9", x"f7", x"09", x"07", x"e0",
    x"f0", x"07", x"14", x"ec", x"d2", x"0e", x"fb", x"fc",
    x"0e", x"19", x"c6", x"e6", x"cb", x"08", x"10", x"bd",
    x"d9", x"15", x"fe", x"05", x"0a", x"d9", x"14", x"17",
    x"e6", x"da", x"02", x"d3", x"15", x"ae", x"fc", x"15",
    x"0e", x"d2", x"dc", x"fa", x"fd", x"01", x"09", x"0a",
    x"fd", x"12", x"fb", x"0b", x"ce", x"0b", x"f9", x"11",
    x"c3", x"09", x"d4", x"09", x"f1", x"17", x"ef", x"d1",
    x"01", x"01", x"cc", x"c5", x"d6", x"d8", x"fc", x"f8",
    x"d6", x"16", x"f5", x"ee", x"02", x"d6", x"10", x"16",
    x"1a", x"0d", x"da", x"fd", x"d3", x"f8", x"f7", x"da",
    x"0f", x"ff", x"fa", x"11", x"0f", x"f4", x"ed", x"fb",
    x"ef", x"07", x"15", x"0d", x"cf", x"13", x"db", x"c8",
    x"f6", x"fd", x"e3", x"c9", x"d0", x"0e", x"fc", x"0c",
    x"10", x"11", x"05", x"e3", x"16", x"d8", x"0d", x"c5",
    x"0b", x"d1", x"e2", x"11", x"cd", x"d7", x"09", x"b4",
    x"13", x"c7", x"0c", x"0a", x"09", x"fe", x"03", x"e0",
    x"0b", x"f6", x"16", x"0b", x"df", x"0e", x"04", x"01",
    x"df", x"13", x"bf", x"d6", x"d7", x"09", x"fb", x"01",
    x"f9", x"cb", x"07", x"fa", x"f9", x"cc", x"d3", x"0b",
    x"cb", x"11", x"fc", x"c6", x"d3", x"00", x"06", x"da",
    x"15", x"11", x"ab", x"06", x"f6", x"fb", x"f1", x"b0",
    x"00", x"16", x"12", x"ff", x"07", x"04", x"f3", x"e0",
    x"ee", x"10", x"c7", x"cf", x"06", x"d5", x"e6", x"0c",
    x"05", x"07", x"9c", x"ba", x"e2", x"e3", x"12", x"07",
    x"12", x"d7", x"0f", x"09", x"ff", x"dc", x"bf", x"d2",
    x"f1", x"0e", x"d6", x"aa", x"f0", x"fe", x"fd", x"ef",
    x"17", x"fa", x"fd", x"06", x"0c", x"05", x"e8", x"f3",
    x"b6", x"ee", x"c6", x"0c", x"c5", x"e2", x"e5", x"da",
    x"ff", x"07", x"0b", x"03", x"e6", x"14", x"00", x"0d",
    x"12", x"c3", x"f9", x"0a", x"de", x"0b", x"15", x"cc",
    x"0f", x"05", x"07", x"19", x"b3", x"1f", x"dd", x"eb",
    x"de", x"c6", x"cd", x"db", x"ff", x"01", x"fb", x"d7",
    x"0b", x"fa", x"0f", x"12", x"0f", x"d5", x"f4", x"f8",
    x"03", x"00", x"09", x"d5", x"ed", x"0a", x"b1", x"03",
    x"ab", x"eb", x"05", x"fb", x"05", x"d8", x"18", x"08",
    x"e1", x"f3", x"01", x"d9", x"08", x"02", x"02", x"33",
    x"dd", x"09", x"0b", x"06", x"05", x"f5", x"0e", x"08",
    x"fa", x"ca", x"f9", x"df", x"e4", x"eb", x"b8", x"16",
    x"d5", x"ca", x"08", x"09", x"fb", x"06", x"10", x"0e",
    x"00", x"05", x"10", x"11", x"0d", x"ff", x"c8", x"04",
    x"f1", x"b9", x"f3", x"1b", x"03", x"0b", x"0f", x"d0",
    x"13", x"cc", x"0d", x"07", x"09", x"ff", x"01", x"d3",
    x"cb", x"f7", x"d6", x"cf", x"f8", x"f7", x"fc", x"f2",
    x"06", x"fd", x"ea", x"c1", x"0d", x"d3", x"0f", x"18",
    x"f7", x"c7", x"06", x"11", x"f6", x"b8", x"f8", x"08",
    x"c9", x"09", x"f7", x"0d", x"19", x"14", x"df", x"f2",
    x"e6", x"dc", x"ce", x"f8", x"0c", x"c1", x"0d", x"09",
    x"ed", x"dd", x"1b", x"09", x"fe", x"13", x"fa", x"1e",
    x"d8", x"f9", x"cc", x"1c", x"e9", x"08", x"01", x"fa",
    x"10", x"15", x"09", x"0f", x"f7", x"b7", x"e2", x"f7",
    x"0e", x"15", x"02", x"fe", x"fb", x"e4", x"de", x"f6",
    x"0d", x"ee", x"07", x"0d", x"d7", x"dc", x"01", x"10",
    x"10", x"ea", x"ff", x"ff", x"f1", x"04", x"17", x"08",
    x"f7", x"12", x"0a", x"fd", x"de", x"f2", x"c6", x"f1",
    x"ed", x"10", x"0c", x"f2", x"05", x"12", x"fe", x"0a",
    x"02", x"0a", x"0a", x"0c", x"c7", x"da", x"db", x"01",
    x"c1", x"0f", x"0f", x"e6", x"06", x"d4", x"db", x"f1",
    x"dd", x"10", x"d6", x"d7", x"0a", x"04", x"04", x"13",
    x"10", x"ef", x"eb", x"d8", x"0e", x"bc", x"d7", x"f9",
    x"e1", x"e2", x"fb", x"08", x"e1", x"ff", x"c4", x"12",
    x"00", x"0d", x"04", x"14", x"9c", x"11", x"00", x"ce",
    x"0f", x"01", x"f6", x"05", x"f2", x"e3", x"09", x"f8",
    x"08", x"db", x"06", x"d7", x"10", x"de", x"e7", x"03",
    x"f1", x"0d", x"e1", x"02", x"00", x"fb", x"02", x"eb",
    x"10", x"f7", x"d4", x"d8", x"c9", x"10", x"f7", x"08",
    x"ea", x"e8", x"0c", x"d5", x"1a", x"0a", x"ff", x"db",
    x"0f", x"f0", x"07", x"06", x"01", x"dd", x"f1", x"e4",
    x"de", x"ee", x"01", x"05", x"ca", x"e2", x"fc", x"cf",
    x"f3", x"d4", x"01", x"fb", x"fb", x"fe", x"eb", x"0d",
    x"f0", x"f5", x"d0", x"cb", x"c1", x"d7", x"c2", x"f5",
    x"e9", x"cd", x"0c", x"02", x"ee", x"de", x"de", x"08",
    x"fd", x"04", x"11", x"0a", x"18", x"00", x"da", x"f9",
    x"06", x"00", x"f2", x"de", x"01", x"0b", x"12", x"e8",
    x"d8", x"d6", x"ef", x"06", x"0a", x"06", x"03", x"14",
    x"c6", x"f1", x"e7", x"08", x"07", x"c0", x"be", x"f5",
    x"f0", x"e3", x"13", x"04", x"12", x"16", x"00", x"13",
    x"fb", x"00", x"d8", x"f3", x"cb", x"cc", x"ee", x"0d",
    x"0b", x"0f", x"0a", x"e5", x"e3", x"15", x"e0", x"0c",
    x"10", x"0a", x"04", x"05", x"0f", x"dc", x"f5", x"09",
    x"d4", x"0c", x"17", x"0b", x"0a", x"e4", x"f8", x"fa",
    x"ef", x"f9", x"ed", x"14", x"d0", x"f8", x"ff", x"fb",
    x"11", x"11", x"dd", x"ed", x"e0", x"09", x"18", x"de",
    x"c6", x"10", x"fa", x"f8", x"fd", x"ee", x"e3", x"10",
    x"e6", x"19", x"01", x"0a", x"1c", x"b6", x"ff", x"12"
  );

  type fc2_bias_10_t is array (0 to 9) of std_logic_vector(7 downto 0);
  constant fc2_bias : fc2_bias_10_t := (
    x"c1", x"2e", x"1e", x"f8", x"15", x"31", x"cf", x"ea",
    x"0e", x"f7"
  );

  type fc2_activation_post_process_eps_1_t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant fc2_activation_post_process_eps : fc2_activation_post_process_eps_1_t := (
    x"00"
  );

  type fc2_activation_post_process_min_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant fc2_activation_post_process_min_val : fc2_activation_post_process_min_val__t := (
    x"83"
  );

  type fc2_activation_post_process_max_val__t is array (0 to 0) of std_logic_vector(7 downto 0);
  constant fc2_activation_post_process_max_val : fc2_activation_post_process_max_val__t := (
    x"57"
  );

end package weights_pkg;
